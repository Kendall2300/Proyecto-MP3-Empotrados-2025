// MP3_PC.v

// Generated using ACDS version 18.0 614

`timescale 1 ps / 1 ps
module MP3_PC (
		input  wire [3:0]  buttons_export_export, // buttons_export.export
		input  wire        clk_clk,               //            clk.clk
		output wire        pll_vga_locked_export, // pll_vga_locked.export
		input  wire        reset_reset_n,         //          reset.reset_n
		output wire [27:0] seven_seg_export,      //      seven_seg.export
		input  wire [2:0]  switchs_export,        //        switchs.export
		output wire        vga_controller_CLK,    // vga_controller.CLK
		output wire        vga_controller_HS,     //               .HS
		output wire        vga_controller_VS,     //               .VS
		output wire        vga_controller_BLANK,  //               .BLANK
		output wire        vga_controller_SYNC,   //               .SYNC
		output wire [7:0]  vga_controller_R,      //               .R
		output wire [7:0]  vga_controller_G,      //               .G
		output wire [7:0]  vga_controller_B       //               .B
	);

	wire         vga_buffer_avalon_char_source_valid;                               // VGA_BUFFER:stream_valid -> VGA_CONTROLLER:valid
	wire  [29:0] vga_buffer_avalon_char_source_data;                                // VGA_BUFFER:stream_data -> VGA_CONTROLLER:data
	wire         vga_buffer_avalon_char_source_ready;                               // VGA_CONTROLLER:ready -> VGA_BUFFER:stream_ready
	wire         vga_buffer_avalon_char_source_startofpacket;                       // VGA_BUFFER:stream_startofpacket -> VGA_CONTROLLER:startofpacket
	wire         vga_buffer_avalon_char_source_endofpacket;                         // VGA_BUFFER:stream_endofpacket -> VGA_CONTROLLER:endofpacket
	wire         pll_vga_outclk0_clk;                                               // PLL_VGA:outclk_0 -> [VGA_BUFFER:clk, VGA_CONTROLLER:clk, mm_interconnect_0:PLL_VGA_outclk0_clk, rst_controller_001:clk]
	wire  [31:0] niosii_data_master_readdata;                                       // mm_interconnect_0:NIOSII_data_master_readdata -> NIOSII:d_readdata
	wire         niosii_data_master_waitrequest;                                    // mm_interconnect_0:NIOSII_data_master_waitrequest -> NIOSII:d_waitrequest
	wire         niosii_data_master_debugaccess;                                    // NIOSII:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:NIOSII_data_master_debugaccess
	wire  [14:0] niosii_data_master_address;                                        // NIOSII:d_address -> mm_interconnect_0:NIOSII_data_master_address
	wire   [3:0] niosii_data_master_byteenable;                                     // NIOSII:d_byteenable -> mm_interconnect_0:NIOSII_data_master_byteenable
	wire         niosii_data_master_read;                                           // NIOSII:d_read -> mm_interconnect_0:NIOSII_data_master_read
	wire         niosii_data_master_write;                                          // NIOSII:d_write -> mm_interconnect_0:NIOSII_data_master_write
	wire  [31:0] niosii_data_master_writedata;                                      // NIOSII:d_writedata -> mm_interconnect_0:NIOSII_data_master_writedata
	wire  [31:0] niosii_instruction_master_readdata;                                // mm_interconnect_0:NIOSII_instruction_master_readdata -> NIOSII:i_readdata
	wire         niosii_instruction_master_waitrequest;                             // mm_interconnect_0:NIOSII_instruction_master_waitrequest -> NIOSII:i_waitrequest
	wire  [14:0] niosii_instruction_master_address;                                 // NIOSII:i_address -> mm_interconnect_0:NIOSII_instruction_master_address
	wire         niosii_instruction_master_read;                                    // NIOSII:i_read -> mm_interconnect_0:NIOSII_instruction_master_read
	wire         mm_interconnect_0_vga_buffer_avalon_char_buffer_slave_chipselect;  // mm_interconnect_0:VGA_BUFFER_avalon_char_buffer_slave_chipselect -> VGA_BUFFER:buf_chipselect
	wire   [7:0] mm_interconnect_0_vga_buffer_avalon_char_buffer_slave_readdata;    // VGA_BUFFER:buf_readdata -> mm_interconnect_0:VGA_BUFFER_avalon_char_buffer_slave_readdata
	wire         mm_interconnect_0_vga_buffer_avalon_char_buffer_slave_waitrequest; // VGA_BUFFER:buf_waitrequest -> mm_interconnect_0:VGA_BUFFER_avalon_char_buffer_slave_waitrequest
	wire  [12:0] mm_interconnect_0_vga_buffer_avalon_char_buffer_slave_address;     // mm_interconnect_0:VGA_BUFFER_avalon_char_buffer_slave_address -> VGA_BUFFER:buf_address
	wire         mm_interconnect_0_vga_buffer_avalon_char_buffer_slave_read;        // mm_interconnect_0:VGA_BUFFER_avalon_char_buffer_slave_read -> VGA_BUFFER:buf_read
	wire   [0:0] mm_interconnect_0_vga_buffer_avalon_char_buffer_slave_byteenable;  // mm_interconnect_0:VGA_BUFFER_avalon_char_buffer_slave_byteenable -> VGA_BUFFER:buf_byteenable
	wire         mm_interconnect_0_vga_buffer_avalon_char_buffer_slave_write;       // mm_interconnect_0:VGA_BUFFER_avalon_char_buffer_slave_write -> VGA_BUFFER:buf_write
	wire   [7:0] mm_interconnect_0_vga_buffer_avalon_char_buffer_slave_writedata;   // mm_interconnect_0:VGA_BUFFER_avalon_char_buffer_slave_writedata -> VGA_BUFFER:buf_writedata
	wire         mm_interconnect_0_vga_buffer_avalon_char_control_slave_chipselect; // mm_interconnect_0:VGA_BUFFER_avalon_char_control_slave_chipselect -> VGA_BUFFER:ctrl_chipselect
	wire  [31:0] mm_interconnect_0_vga_buffer_avalon_char_control_slave_readdata;   // VGA_BUFFER:ctrl_readdata -> mm_interconnect_0:VGA_BUFFER_avalon_char_control_slave_readdata
	wire   [0:0] mm_interconnect_0_vga_buffer_avalon_char_control_slave_address;    // mm_interconnect_0:VGA_BUFFER_avalon_char_control_slave_address -> VGA_BUFFER:ctrl_address
	wire         mm_interconnect_0_vga_buffer_avalon_char_control_slave_read;       // mm_interconnect_0:VGA_BUFFER_avalon_char_control_slave_read -> VGA_BUFFER:ctrl_read
	wire   [3:0] mm_interconnect_0_vga_buffer_avalon_char_control_slave_byteenable; // mm_interconnect_0:VGA_BUFFER_avalon_char_control_slave_byteenable -> VGA_BUFFER:ctrl_byteenable
	wire         mm_interconnect_0_vga_buffer_avalon_char_control_slave_write;      // mm_interconnect_0:VGA_BUFFER_avalon_char_control_slave_write -> VGA_BUFFER:ctrl_write
	wire  [31:0] mm_interconnect_0_vga_buffer_avalon_char_control_slave_writedata;  // mm_interconnect_0:VGA_BUFFER_avalon_char_control_slave_writedata -> VGA_BUFFER:ctrl_writedata
	wire         mm_interconnect_0_uart_avalon_jtag_slave_chipselect;               // mm_interconnect_0:UART_avalon_jtag_slave_chipselect -> UART:av_chipselect
	wire  [31:0] mm_interconnect_0_uart_avalon_jtag_slave_readdata;                 // UART:av_readdata -> mm_interconnect_0:UART_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_uart_avalon_jtag_slave_waitrequest;              // UART:av_waitrequest -> mm_interconnect_0:UART_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_uart_avalon_jtag_slave_address;                  // mm_interconnect_0:UART_avalon_jtag_slave_address -> UART:av_address
	wire         mm_interconnect_0_uart_avalon_jtag_slave_read;                     // mm_interconnect_0:UART_avalon_jtag_slave_read -> UART:av_read_n
	wire         mm_interconnect_0_uart_avalon_jtag_slave_write;                    // mm_interconnect_0:UART_avalon_jtag_slave_write -> UART:av_write_n
	wire  [31:0] mm_interconnect_0_uart_avalon_jtag_slave_writedata;                // mm_interconnect_0:UART_avalon_jtag_slave_writedata -> UART:av_writedata
	wire  [31:0] mm_interconnect_0_niosii_debug_mem_slave_readdata;                 // NIOSII:debug_mem_slave_readdata -> mm_interconnect_0:NIOSII_debug_mem_slave_readdata
	wire         mm_interconnect_0_niosii_debug_mem_slave_waitrequest;              // NIOSII:debug_mem_slave_waitrequest -> mm_interconnect_0:NIOSII_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_niosii_debug_mem_slave_debugaccess;              // mm_interconnect_0:NIOSII_debug_mem_slave_debugaccess -> NIOSII:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_niosii_debug_mem_slave_address;                  // mm_interconnect_0:NIOSII_debug_mem_slave_address -> NIOSII:debug_mem_slave_address
	wire         mm_interconnect_0_niosii_debug_mem_slave_read;                     // mm_interconnect_0:NIOSII_debug_mem_slave_read -> NIOSII:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_niosii_debug_mem_slave_byteenable;               // mm_interconnect_0:NIOSII_debug_mem_slave_byteenable -> NIOSII:debug_mem_slave_byteenable
	wire         mm_interconnect_0_niosii_debug_mem_slave_write;                    // mm_interconnect_0:NIOSII_debug_mem_slave_write -> NIOSII:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_niosii_debug_mem_slave_writedata;                // mm_interconnect_0:NIOSII_debug_mem_slave_writedata -> NIOSII:debug_mem_slave_writedata
	wire         mm_interconnect_0_timer_1s_s1_chipselect;                          // mm_interconnect_0:TIMER_1s_s1_chipselect -> TIMER_1s:chipselect
	wire  [15:0] mm_interconnect_0_timer_1s_s1_readdata;                            // TIMER_1s:readdata -> mm_interconnect_0:TIMER_1s_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_1s_s1_address;                             // mm_interconnect_0:TIMER_1s_s1_address -> TIMER_1s:address
	wire         mm_interconnect_0_timer_1s_s1_write;                               // mm_interconnect_0:TIMER_1s_s1_write -> TIMER_1s:write_n
	wire  [15:0] mm_interconnect_0_timer_1s_s1_writedata;                           // mm_interconnect_0:TIMER_1s_s1_writedata -> TIMER_1s:writedata
	wire         mm_interconnect_0_reg_7seg_s1_chipselect;                          // mm_interconnect_0:REG_7SEG_s1_chipselect -> REG_7SEG:chipselect
	wire  [31:0] mm_interconnect_0_reg_7seg_s1_readdata;                            // REG_7SEG:readdata -> mm_interconnect_0:REG_7SEG_s1_readdata
	wire   [1:0] mm_interconnect_0_reg_7seg_s1_address;                             // mm_interconnect_0:REG_7SEG_s1_address -> REG_7SEG:address
	wire         mm_interconnect_0_reg_7seg_s1_write;                               // mm_interconnect_0:REG_7SEG_s1_write -> REG_7SEG:write_n
	wire  [31:0] mm_interconnect_0_reg_7seg_s1_writedata;                           // mm_interconnect_0:REG_7SEG_s1_writedata -> REG_7SEG:writedata
	wire  [31:0] mm_interconnect_0_reg_switch_s1_readdata;                          // REG_SWITCH:readdata -> mm_interconnect_0:REG_SWITCH_s1_readdata
	wire   [1:0] mm_interconnect_0_reg_switch_s1_address;                           // mm_interconnect_0:REG_SWITCH_s1_address -> REG_SWITCH:address
	wire         mm_interconnect_0_reg_button_s1_chipselect;                        // mm_interconnect_0:REG_BUTTON_s1_chipselect -> REG_BUTTON:chipselect
	wire  [31:0] mm_interconnect_0_reg_button_s1_readdata;                          // REG_BUTTON:readdata -> mm_interconnect_0:REG_BUTTON_s1_readdata
	wire   [1:0] mm_interconnect_0_reg_button_s1_address;                           // mm_interconnect_0:REG_BUTTON_s1_address -> REG_BUTTON:address
	wire         mm_interconnect_0_reg_button_s1_write;                             // mm_interconnect_0:REG_BUTTON_s1_write -> REG_BUTTON:write_n
	wire  [31:0] mm_interconnect_0_reg_button_s1_writedata;                         // mm_interconnect_0:REG_BUTTON_s1_writedata -> REG_BUTTON:writedata
	wire         mm_interconnect_0_ram_s1_chipselect;                               // mm_interconnect_0:RAM_s1_chipselect -> RAM:chipselect
	wire  [31:0] mm_interconnect_0_ram_s1_readdata;                                 // RAM:readdata -> mm_interconnect_0:RAM_s1_readdata
	wire  [11:0] mm_interconnect_0_ram_s1_address;                                  // mm_interconnect_0:RAM_s1_address -> RAM:address
	wire   [3:0] mm_interconnect_0_ram_s1_byteenable;                               // mm_interconnect_0:RAM_s1_byteenable -> RAM:byteenable
	wire         mm_interconnect_0_ram_s1_write;                                    // mm_interconnect_0:RAM_s1_write -> RAM:write
	wire  [31:0] mm_interconnect_0_ram_s1_writedata;                                // mm_interconnect_0:RAM_s1_writedata -> RAM:writedata
	wire         mm_interconnect_0_ram_s1_clken;                                    // mm_interconnect_0:RAM_s1_clken -> RAM:clken
	wire         irq_mapper_receiver0_irq;                                          // TIMER_1s:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                          // REG_BUTTON:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                          // UART:av_irq -> irq_mapper:receiver2_irq
	wire  [31:0] niosii_irq_irq;                                                    // irq_mapper:sender_irq -> NIOSII:irq
	wire         rst_controller_reset_out_reset;                                    // rst_controller:reset_out -> [NIOSII:reset_n, RAM:reset, REG_7SEG:reset_n, REG_BUTTON:reset_n, REG_SWITCH:reset_n, TIMER_1s:reset_n, UART:rst_n, irq_mapper:reset, mm_interconnect_0:NIOSII_reset_reset_bridge_in_reset_reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                                // rst_controller:reset_req -> [NIOSII:reset_req, RAM:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_001_reset_out_reset;                                // rst_controller_001:reset_out -> [VGA_BUFFER:reset, VGA_CONTROLLER:reset, mm_interconnect_0:VGA_BUFFER_reset_reset_bridge_in_reset_reset]

	MP3_PC_NIOSII niosii (
		.clk                                 (clk_clk),                                              //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                      //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                   //                          .reset_req
		.d_address                           (niosii_data_master_address),                           //               data_master.address
		.d_byteenable                        (niosii_data_master_byteenable),                        //                          .byteenable
		.d_read                              (niosii_data_master_read),                              //                          .read
		.d_readdata                          (niosii_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (niosii_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (niosii_data_master_write),                             //                          .write
		.d_writedata                         (niosii_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (niosii_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (niosii_instruction_master_address),                    //        instruction_master.address
		.i_read                              (niosii_instruction_master_read),                       //                          .read
		.i_readdata                          (niosii_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (niosii_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (niosii_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_niosii_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_niosii_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_niosii_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_niosii_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_niosii_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_niosii_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_niosii_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_niosii_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                      // custom_instruction_master.readra
	);

	MP3_PC_PLL_VGA pll_vga (
		.refclk   (clk_clk),               //  refclk.clk
		.rst      (~reset_reset_n),        //   reset.reset
		.outclk_0 (pll_vga_outclk0_clk),   // outclk0.clk
		.locked   (pll_vga_locked_export)  //  locked.export
	);

	MP3_PC_RAM ram (
		.clk        (clk_clk),                             //   clk1.clk
		.address    (mm_interconnect_0_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),      // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),  //       .reset_req
		.freeze     (1'b0)                                 // (terminated)
	);

	MP3_PC_REG_7SEG reg_7seg (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_reg_7seg_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_reg_7seg_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_reg_7seg_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_reg_7seg_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_reg_7seg_s1_readdata),   //                    .readdata
		.out_port   (seven_seg_export)                          // external_connection.export
	);

	MP3_PC_REG_BUTTON reg_button (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_reg_button_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_reg_button_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_reg_button_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_reg_button_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_reg_button_s1_readdata),   //                    .readdata
		.in_port    (buttons_export_export),                      // external_connection.export
		.irq        (irq_mapper_receiver1_irq)                    //                 irq.irq
	);

	MP3_PC_REG_SWITCH reg_switch (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address  (mm_interconnect_0_reg_switch_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_reg_switch_s1_readdata), //                    .readdata
		.in_port  (switchs_export)                            // external_connection.export
	);

	MP3_PC_TIMER_1s timer_1s (
		.clk        (clk_clk),                                  //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          // reset.reset_n
		.address    (mm_interconnect_0_timer_1s_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_1s_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_1s_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_1s_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_1s_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)                  //   irq.irq
	);

	MP3_PC_UART uart (
		.clk            (clk_clk),                                              //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                      //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver2_irq)                              //               irq.irq
	);

	MP3_PC_VGA_BUFFER vga_buffer (
		.clk                  (pll_vga_outclk0_clk),                                               //                       clk.clk
		.reset                (rst_controller_001_reset_out_reset),                                //                     reset.reset
		.ctrl_address         (mm_interconnect_0_vga_buffer_avalon_char_control_slave_address),    // avalon_char_control_slave.address
		.ctrl_byteenable      (mm_interconnect_0_vga_buffer_avalon_char_control_slave_byteenable), //                          .byteenable
		.ctrl_chipselect      (mm_interconnect_0_vga_buffer_avalon_char_control_slave_chipselect), //                          .chipselect
		.ctrl_read            (mm_interconnect_0_vga_buffer_avalon_char_control_slave_read),       //                          .read
		.ctrl_write           (mm_interconnect_0_vga_buffer_avalon_char_control_slave_write),      //                          .write
		.ctrl_writedata       (mm_interconnect_0_vga_buffer_avalon_char_control_slave_writedata),  //                          .writedata
		.ctrl_readdata        (mm_interconnect_0_vga_buffer_avalon_char_control_slave_readdata),   //                          .readdata
		.buf_byteenable       (mm_interconnect_0_vga_buffer_avalon_char_buffer_slave_byteenable),  //  avalon_char_buffer_slave.byteenable
		.buf_chipselect       (mm_interconnect_0_vga_buffer_avalon_char_buffer_slave_chipselect),  //                          .chipselect
		.buf_read             (mm_interconnect_0_vga_buffer_avalon_char_buffer_slave_read),        //                          .read
		.buf_write            (mm_interconnect_0_vga_buffer_avalon_char_buffer_slave_write),       //                          .write
		.buf_writedata        (mm_interconnect_0_vga_buffer_avalon_char_buffer_slave_writedata),   //                          .writedata
		.buf_readdata         (mm_interconnect_0_vga_buffer_avalon_char_buffer_slave_readdata),    //                          .readdata
		.buf_waitrequest      (mm_interconnect_0_vga_buffer_avalon_char_buffer_slave_waitrequest), //                          .waitrequest
		.buf_address          (mm_interconnect_0_vga_buffer_avalon_char_buffer_slave_address),     //                          .address
		.stream_ready         (vga_buffer_avalon_char_source_ready),                               //        avalon_char_source.ready
		.stream_startofpacket (vga_buffer_avalon_char_source_startofpacket),                       //                          .startofpacket
		.stream_endofpacket   (vga_buffer_avalon_char_source_endofpacket),                         //                          .endofpacket
		.stream_valid         (vga_buffer_avalon_char_source_valid),                               //                          .valid
		.stream_data          (vga_buffer_avalon_char_source_data)                                 //                          .data
	);

	MP3_PC_VGA_CONTROLLER vga_controller (
		.clk           (pll_vga_outclk0_clk),                         //                clk.clk
		.reset         (rst_controller_001_reset_out_reset),          //              reset.reset
		.data          (vga_buffer_avalon_char_source_data),          //    avalon_vga_sink.data
		.startofpacket (vga_buffer_avalon_char_source_startofpacket), //                   .startofpacket
		.endofpacket   (vga_buffer_avalon_char_source_endofpacket),   //                   .endofpacket
		.valid         (vga_buffer_avalon_char_source_valid),         //                   .valid
		.ready         (vga_buffer_avalon_char_source_ready),         //                   .ready
		.VGA_CLK       (vga_controller_CLK),                          // external_interface.export
		.VGA_HS        (vga_controller_HS),                           //                   .export
		.VGA_VS        (vga_controller_VS),                           //                   .export
		.VGA_BLANK     (vga_controller_BLANK),                        //                   .export
		.VGA_SYNC      (vga_controller_SYNC),                         //                   .export
		.VGA_R         (vga_controller_R),                            //                   .export
		.VGA_G         (vga_controller_G),                            //                   .export
		.VGA_B         (vga_controller_B)                             //                   .export
	);

	MP3_PC_mm_interconnect_0 mm_interconnect_0 (
		.CLK_clk_clk                                     (clk_clk),                                                           //                                CLK_clk.clk
		.PLL_VGA_outclk0_clk                             (pll_vga_outclk0_clk),                                               //                        PLL_VGA_outclk0.clk
		.NIOSII_reset_reset_bridge_in_reset_reset        (rst_controller_reset_out_reset),                                    //     NIOSII_reset_reset_bridge_in_reset.reset
		.VGA_BUFFER_reset_reset_bridge_in_reset_reset    (rst_controller_001_reset_out_reset),                                // VGA_BUFFER_reset_reset_bridge_in_reset.reset
		.NIOSII_data_master_address                      (niosii_data_master_address),                                        //                     NIOSII_data_master.address
		.NIOSII_data_master_waitrequest                  (niosii_data_master_waitrequest),                                    //                                       .waitrequest
		.NIOSII_data_master_byteenable                   (niosii_data_master_byteenable),                                     //                                       .byteenable
		.NIOSII_data_master_read                         (niosii_data_master_read),                                           //                                       .read
		.NIOSII_data_master_readdata                     (niosii_data_master_readdata),                                       //                                       .readdata
		.NIOSII_data_master_write                        (niosii_data_master_write),                                          //                                       .write
		.NIOSII_data_master_writedata                    (niosii_data_master_writedata),                                      //                                       .writedata
		.NIOSII_data_master_debugaccess                  (niosii_data_master_debugaccess),                                    //                                       .debugaccess
		.NIOSII_instruction_master_address               (niosii_instruction_master_address),                                 //              NIOSII_instruction_master.address
		.NIOSII_instruction_master_waitrequest           (niosii_instruction_master_waitrequest),                             //                                       .waitrequest
		.NIOSII_instruction_master_read                  (niosii_instruction_master_read),                                    //                                       .read
		.NIOSII_instruction_master_readdata              (niosii_instruction_master_readdata),                                //                                       .readdata
		.NIOSII_debug_mem_slave_address                  (mm_interconnect_0_niosii_debug_mem_slave_address),                  //                 NIOSII_debug_mem_slave.address
		.NIOSII_debug_mem_slave_write                    (mm_interconnect_0_niosii_debug_mem_slave_write),                    //                                       .write
		.NIOSII_debug_mem_slave_read                     (mm_interconnect_0_niosii_debug_mem_slave_read),                     //                                       .read
		.NIOSII_debug_mem_slave_readdata                 (mm_interconnect_0_niosii_debug_mem_slave_readdata),                 //                                       .readdata
		.NIOSII_debug_mem_slave_writedata                (mm_interconnect_0_niosii_debug_mem_slave_writedata),                //                                       .writedata
		.NIOSII_debug_mem_slave_byteenable               (mm_interconnect_0_niosii_debug_mem_slave_byteenable),               //                                       .byteenable
		.NIOSII_debug_mem_slave_waitrequest              (mm_interconnect_0_niosii_debug_mem_slave_waitrequest),              //                                       .waitrequest
		.NIOSII_debug_mem_slave_debugaccess              (mm_interconnect_0_niosii_debug_mem_slave_debugaccess),              //                                       .debugaccess
		.RAM_s1_address                                  (mm_interconnect_0_ram_s1_address),                                  //                                 RAM_s1.address
		.RAM_s1_write                                    (mm_interconnect_0_ram_s1_write),                                    //                                       .write
		.RAM_s1_readdata                                 (mm_interconnect_0_ram_s1_readdata),                                 //                                       .readdata
		.RAM_s1_writedata                                (mm_interconnect_0_ram_s1_writedata),                                //                                       .writedata
		.RAM_s1_byteenable                               (mm_interconnect_0_ram_s1_byteenable),                               //                                       .byteenable
		.RAM_s1_chipselect                               (mm_interconnect_0_ram_s1_chipselect),                               //                                       .chipselect
		.RAM_s1_clken                                    (mm_interconnect_0_ram_s1_clken),                                    //                                       .clken
		.REG_7SEG_s1_address                             (mm_interconnect_0_reg_7seg_s1_address),                             //                            REG_7SEG_s1.address
		.REG_7SEG_s1_write                               (mm_interconnect_0_reg_7seg_s1_write),                               //                                       .write
		.REG_7SEG_s1_readdata                            (mm_interconnect_0_reg_7seg_s1_readdata),                            //                                       .readdata
		.REG_7SEG_s1_writedata                           (mm_interconnect_0_reg_7seg_s1_writedata),                           //                                       .writedata
		.REG_7SEG_s1_chipselect                          (mm_interconnect_0_reg_7seg_s1_chipselect),                          //                                       .chipselect
		.REG_BUTTON_s1_address                           (mm_interconnect_0_reg_button_s1_address),                           //                          REG_BUTTON_s1.address
		.REG_BUTTON_s1_write                             (mm_interconnect_0_reg_button_s1_write),                             //                                       .write
		.REG_BUTTON_s1_readdata                          (mm_interconnect_0_reg_button_s1_readdata),                          //                                       .readdata
		.REG_BUTTON_s1_writedata                         (mm_interconnect_0_reg_button_s1_writedata),                         //                                       .writedata
		.REG_BUTTON_s1_chipselect                        (mm_interconnect_0_reg_button_s1_chipselect),                        //                                       .chipselect
		.REG_SWITCH_s1_address                           (mm_interconnect_0_reg_switch_s1_address),                           //                          REG_SWITCH_s1.address
		.REG_SWITCH_s1_readdata                          (mm_interconnect_0_reg_switch_s1_readdata),                          //                                       .readdata
		.TIMER_1s_s1_address                             (mm_interconnect_0_timer_1s_s1_address),                             //                            TIMER_1s_s1.address
		.TIMER_1s_s1_write                               (mm_interconnect_0_timer_1s_s1_write),                               //                                       .write
		.TIMER_1s_s1_readdata                            (mm_interconnect_0_timer_1s_s1_readdata),                            //                                       .readdata
		.TIMER_1s_s1_writedata                           (mm_interconnect_0_timer_1s_s1_writedata),                           //                                       .writedata
		.TIMER_1s_s1_chipselect                          (mm_interconnect_0_timer_1s_s1_chipselect),                          //                                       .chipselect
		.UART_avalon_jtag_slave_address                  (mm_interconnect_0_uart_avalon_jtag_slave_address),                  //                 UART_avalon_jtag_slave.address
		.UART_avalon_jtag_slave_write                    (mm_interconnect_0_uart_avalon_jtag_slave_write),                    //                                       .write
		.UART_avalon_jtag_slave_read                     (mm_interconnect_0_uart_avalon_jtag_slave_read),                     //                                       .read
		.UART_avalon_jtag_slave_readdata                 (mm_interconnect_0_uart_avalon_jtag_slave_readdata),                 //                                       .readdata
		.UART_avalon_jtag_slave_writedata                (mm_interconnect_0_uart_avalon_jtag_slave_writedata),                //                                       .writedata
		.UART_avalon_jtag_slave_waitrequest              (mm_interconnect_0_uart_avalon_jtag_slave_waitrequest),              //                                       .waitrequest
		.UART_avalon_jtag_slave_chipselect               (mm_interconnect_0_uart_avalon_jtag_slave_chipselect),               //                                       .chipselect
		.VGA_BUFFER_avalon_char_buffer_slave_address     (mm_interconnect_0_vga_buffer_avalon_char_buffer_slave_address),     //    VGA_BUFFER_avalon_char_buffer_slave.address
		.VGA_BUFFER_avalon_char_buffer_slave_write       (mm_interconnect_0_vga_buffer_avalon_char_buffer_slave_write),       //                                       .write
		.VGA_BUFFER_avalon_char_buffer_slave_read        (mm_interconnect_0_vga_buffer_avalon_char_buffer_slave_read),        //                                       .read
		.VGA_BUFFER_avalon_char_buffer_slave_readdata    (mm_interconnect_0_vga_buffer_avalon_char_buffer_slave_readdata),    //                                       .readdata
		.VGA_BUFFER_avalon_char_buffer_slave_writedata   (mm_interconnect_0_vga_buffer_avalon_char_buffer_slave_writedata),   //                                       .writedata
		.VGA_BUFFER_avalon_char_buffer_slave_byteenable  (mm_interconnect_0_vga_buffer_avalon_char_buffer_slave_byteenable),  //                                       .byteenable
		.VGA_BUFFER_avalon_char_buffer_slave_waitrequest (mm_interconnect_0_vga_buffer_avalon_char_buffer_slave_waitrequest), //                                       .waitrequest
		.VGA_BUFFER_avalon_char_buffer_slave_chipselect  (mm_interconnect_0_vga_buffer_avalon_char_buffer_slave_chipselect),  //                                       .chipselect
		.VGA_BUFFER_avalon_char_control_slave_address    (mm_interconnect_0_vga_buffer_avalon_char_control_slave_address),    //   VGA_BUFFER_avalon_char_control_slave.address
		.VGA_BUFFER_avalon_char_control_slave_write      (mm_interconnect_0_vga_buffer_avalon_char_control_slave_write),      //                                       .write
		.VGA_BUFFER_avalon_char_control_slave_read       (mm_interconnect_0_vga_buffer_avalon_char_control_slave_read),       //                                       .read
		.VGA_BUFFER_avalon_char_control_slave_readdata   (mm_interconnect_0_vga_buffer_avalon_char_control_slave_readdata),   //                                       .readdata
		.VGA_BUFFER_avalon_char_control_slave_writedata  (mm_interconnect_0_vga_buffer_avalon_char_control_slave_writedata),  //                                       .writedata
		.VGA_BUFFER_avalon_char_control_slave_byteenable (mm_interconnect_0_vga_buffer_avalon_char_control_slave_byteenable), //                                       .byteenable
		.VGA_BUFFER_avalon_char_control_slave_chipselect (mm_interconnect_0_vga_buffer_avalon_char_control_slave_chipselect)  //                                       .chipselect
	);

	MP3_PC_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.sender_irq    (niosii_irq_irq)                  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (pll_vga_outclk0_clk),                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
