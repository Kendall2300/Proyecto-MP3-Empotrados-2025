// MP3_PC.v

// Generated using ACDS version 18.0 614

`timescale 1 ps / 1 ps
module MP3_PC (
		inout  wire        audio_config_SDAT,             //       audio_config.SDAT
		output wire        audio_config_SCLK,             //                   .SCLK
		input  wire        audio_external_BCLK,           //     audio_external.BCLK
		output wire        audio_external_DACDAT,         //                   .DACDAT
		input  wire        audio_external_DACLRCK,        //                   .DACLRCK
		output wire        audio_pll_clk_clk,             //      audio_pll_clk.clk
		input  wire [3:0]  buttons_export_export,         //     buttons_export.export
		input  wire        clk_clk,                       //                clk.clk
		input  wire        hps_h2f_mpu_events_eventi,     // hps_h2f_mpu_events.eventi
		output wire        hps_h2f_mpu_events_evento,     //                   .evento
		output wire [1:0]  hps_h2f_mpu_events_standbywfe, //                   .standbywfe
		output wire [1:0]  hps_h2f_mpu_events_standbywfi, //                   .standbywfi
		inout  wire        hps_io_hps_io_sdio_inst_CMD,   //             hps_io.hps_io_sdio_inst_CMD
		inout  wire        hps_io_hps_io_sdio_inst_D0,    //                   .hps_io_sdio_inst_D0
		inout  wire        hps_io_hps_io_sdio_inst_D1,    //                   .hps_io_sdio_inst_D1
		output wire        hps_io_hps_io_sdio_inst_CLK,   //                   .hps_io_sdio_inst_CLK
		inout  wire        hps_io_hps_io_sdio_inst_D2,    //                   .hps_io_sdio_inst_D2
		inout  wire        hps_io_hps_io_sdio_inst_D3,    //                   .hps_io_sdio_inst_D3
		output wire [12:0] memory_mem_a,                  //             memory.mem_a
		output wire [2:0]  memory_mem_ba,                 //                   .mem_ba
		output wire        memory_mem_ck,                 //                   .mem_ck
		output wire        memory_mem_ck_n,               //                   .mem_ck_n
		output wire        memory_mem_cke,                //                   .mem_cke
		output wire        memory_mem_cs_n,               //                   .mem_cs_n
		output wire        memory_mem_ras_n,              //                   .mem_ras_n
		output wire        memory_mem_cas_n,              //                   .mem_cas_n
		output wire        memory_mem_we_n,               //                   .mem_we_n
		output wire        memory_mem_reset_n,            //                   .mem_reset_n
		inout  wire [7:0]  memory_mem_dq,                 //                   .mem_dq
		inout  wire        memory_mem_dqs,                //                   .mem_dqs
		inout  wire        memory_mem_dqs_n,              //                   .mem_dqs_n
		output wire        memory_mem_odt,                //                   .mem_odt
		output wire        memory_mem_dm,                 //                   .mem_dm
		input  wire        memory_oct_rzqin,              //                   .oct_rzqin
		output wire        pll_vga_locked_export,         //     pll_vga_locked.export
		output wire [27:0] seven_seg_export,              //          seven_seg.export
		input  wire [2:0]  switchs_export,                //            switchs.export
		output wire        vga_controller_CLK,            //     vga_controller.CLK
		output wire        vga_controller_HS,             //                   .HS
		output wire        vga_controller_VS,             //                   .VS
		output wire        vga_controller_BLANK,          //                   .BLANK
		output wire        vga_controller_SYNC,           //                   .SYNC
		output wire [7:0]  vga_controller_R,              //                   .R
		output wire [7:0]  vga_controller_G,              //                   .G
		output wire [7:0]  vga_controller_B               //                   .B
	);

	wire         vga_buffer_avalon_char_source_valid;                               // VGA_BUFFER:stream_valid -> VGA_CONTROLLER:valid
	wire  [29:0] vga_buffer_avalon_char_source_data;                                // VGA_BUFFER:stream_data -> VGA_CONTROLLER:data
	wire         vga_buffer_avalon_char_source_ready;                               // VGA_CONTROLLER:ready -> VGA_BUFFER:stream_ready
	wire         vga_buffer_avalon_char_source_startofpacket;                       // VGA_BUFFER:stream_startofpacket -> VGA_CONTROLLER:startofpacket
	wire         vga_buffer_avalon_char_source_endofpacket;                         // VGA_BUFFER:stream_endofpacket -> VGA_CONTROLLER:endofpacket
	wire         pll_vga_outclk0_clk;                                               // PLL_VGA:outclk_0 -> [VGA_BUFFER:clk, VGA_CONTROLLER:clk, mm_interconnect_0:PLL_VGA_outclk0_clk, rst_controller_002:clk]
	wire         hps_h2f_reset_reset;                                               // HPS:h2f_rst_n -> [AudioPLL:ref_reset_reset, PLL_VGA:rst, rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0]
	wire  [31:0] niosii_data_master_readdata;                                       // mm_interconnect_0:NIOSII_data_master_readdata -> NIOSII:d_readdata
	wire         niosii_data_master_waitrequest;                                    // mm_interconnect_0:NIOSII_data_master_waitrequest -> NIOSII:d_waitrequest
	wire         niosii_data_master_debugaccess;                                    // NIOSII:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:NIOSII_data_master_debugaccess
	wire  [15:0] niosii_data_master_address;                                        // NIOSII:d_address -> mm_interconnect_0:NIOSII_data_master_address
	wire   [3:0] niosii_data_master_byteenable;                                     // NIOSII:d_byteenable -> mm_interconnect_0:NIOSII_data_master_byteenable
	wire         niosii_data_master_read;                                           // NIOSII:d_read -> mm_interconnect_0:NIOSII_data_master_read
	wire         niosii_data_master_write;                                          // NIOSII:d_write -> mm_interconnect_0:NIOSII_data_master_write
	wire  [31:0] niosii_data_master_writedata;                                      // NIOSII:d_writedata -> mm_interconnect_0:NIOSII_data_master_writedata
	wire  [31:0] niosii_instruction_master_readdata;                                // mm_interconnect_0:NIOSII_instruction_master_readdata -> NIOSII:i_readdata
	wire         niosii_instruction_master_waitrequest;                             // mm_interconnect_0:NIOSII_instruction_master_waitrequest -> NIOSII:i_waitrequest
	wire  [14:0] niosii_instruction_master_address;                                 // NIOSII:i_address -> mm_interconnect_0:NIOSII_instruction_master_address
	wire         niosii_instruction_master_read;                                    // NIOSII:i_read -> mm_interconnect_0:NIOSII_instruction_master_read
	wire         mm_interconnect_0_audio_avalon_audio_slave_chipselect;             // mm_interconnect_0:Audio_avalon_audio_slave_chipselect -> Audio:chipselect
	wire  [31:0] mm_interconnect_0_audio_avalon_audio_slave_readdata;               // Audio:readdata -> mm_interconnect_0:Audio_avalon_audio_slave_readdata
	wire   [1:0] mm_interconnect_0_audio_avalon_audio_slave_address;                // mm_interconnect_0:Audio_avalon_audio_slave_address -> Audio:address
	wire         mm_interconnect_0_audio_avalon_audio_slave_read;                   // mm_interconnect_0:Audio_avalon_audio_slave_read -> Audio:read
	wire         mm_interconnect_0_audio_avalon_audio_slave_write;                  // mm_interconnect_0:Audio_avalon_audio_slave_write -> Audio:write
	wire  [31:0] mm_interconnect_0_audio_avalon_audio_slave_writedata;              // mm_interconnect_0:Audio_avalon_audio_slave_writedata -> Audio:writedata
	wire  [31:0] mm_interconnect_0_audioconfig_avalon_av_config_slave_readdata;     // AudioConfig:readdata -> mm_interconnect_0:AudioConfig_avalon_av_config_slave_readdata
	wire         mm_interconnect_0_audioconfig_avalon_av_config_slave_waitrequest;  // AudioConfig:waitrequest -> mm_interconnect_0:AudioConfig_avalon_av_config_slave_waitrequest
	wire   [1:0] mm_interconnect_0_audioconfig_avalon_av_config_slave_address;      // mm_interconnect_0:AudioConfig_avalon_av_config_slave_address -> AudioConfig:address
	wire         mm_interconnect_0_audioconfig_avalon_av_config_slave_read;         // mm_interconnect_0:AudioConfig_avalon_av_config_slave_read -> AudioConfig:read
	wire   [3:0] mm_interconnect_0_audioconfig_avalon_av_config_slave_byteenable;   // mm_interconnect_0:AudioConfig_avalon_av_config_slave_byteenable -> AudioConfig:byteenable
	wire         mm_interconnect_0_audioconfig_avalon_av_config_slave_write;        // mm_interconnect_0:AudioConfig_avalon_av_config_slave_write -> AudioConfig:write
	wire  [31:0] mm_interconnect_0_audioconfig_avalon_av_config_slave_writedata;    // mm_interconnect_0:AudioConfig_avalon_av_config_slave_writedata -> AudioConfig:writedata
	wire         mm_interconnect_0_vga_buffer_avalon_char_buffer_slave_chipselect;  // mm_interconnect_0:VGA_BUFFER_avalon_char_buffer_slave_chipselect -> VGA_BUFFER:buf_chipselect
	wire   [7:0] mm_interconnect_0_vga_buffer_avalon_char_buffer_slave_readdata;    // VGA_BUFFER:buf_readdata -> mm_interconnect_0:VGA_BUFFER_avalon_char_buffer_slave_readdata
	wire         mm_interconnect_0_vga_buffer_avalon_char_buffer_slave_waitrequest; // VGA_BUFFER:buf_waitrequest -> mm_interconnect_0:VGA_BUFFER_avalon_char_buffer_slave_waitrequest
	wire  [12:0] mm_interconnect_0_vga_buffer_avalon_char_buffer_slave_address;     // mm_interconnect_0:VGA_BUFFER_avalon_char_buffer_slave_address -> VGA_BUFFER:buf_address
	wire         mm_interconnect_0_vga_buffer_avalon_char_buffer_slave_read;        // mm_interconnect_0:VGA_BUFFER_avalon_char_buffer_slave_read -> VGA_BUFFER:buf_read
	wire   [0:0] mm_interconnect_0_vga_buffer_avalon_char_buffer_slave_byteenable;  // mm_interconnect_0:VGA_BUFFER_avalon_char_buffer_slave_byteenable -> VGA_BUFFER:buf_byteenable
	wire         mm_interconnect_0_vga_buffer_avalon_char_buffer_slave_write;       // mm_interconnect_0:VGA_BUFFER_avalon_char_buffer_slave_write -> VGA_BUFFER:buf_write
	wire   [7:0] mm_interconnect_0_vga_buffer_avalon_char_buffer_slave_writedata;   // mm_interconnect_0:VGA_BUFFER_avalon_char_buffer_slave_writedata -> VGA_BUFFER:buf_writedata
	wire         mm_interconnect_0_vga_buffer_avalon_char_control_slave_chipselect; // mm_interconnect_0:VGA_BUFFER_avalon_char_control_slave_chipselect -> VGA_BUFFER:ctrl_chipselect
	wire  [31:0] mm_interconnect_0_vga_buffer_avalon_char_control_slave_readdata;   // VGA_BUFFER:ctrl_readdata -> mm_interconnect_0:VGA_BUFFER_avalon_char_control_slave_readdata
	wire   [0:0] mm_interconnect_0_vga_buffer_avalon_char_control_slave_address;    // mm_interconnect_0:VGA_BUFFER_avalon_char_control_slave_address -> VGA_BUFFER:ctrl_address
	wire         mm_interconnect_0_vga_buffer_avalon_char_control_slave_read;       // mm_interconnect_0:VGA_BUFFER_avalon_char_control_slave_read -> VGA_BUFFER:ctrl_read
	wire   [3:0] mm_interconnect_0_vga_buffer_avalon_char_control_slave_byteenable; // mm_interconnect_0:VGA_BUFFER_avalon_char_control_slave_byteenable -> VGA_BUFFER:ctrl_byteenable
	wire         mm_interconnect_0_vga_buffer_avalon_char_control_slave_write;      // mm_interconnect_0:VGA_BUFFER_avalon_char_control_slave_write -> VGA_BUFFER:ctrl_write
	wire  [31:0] mm_interconnect_0_vga_buffer_avalon_char_control_slave_writedata;  // mm_interconnect_0:VGA_BUFFER_avalon_char_control_slave_writedata -> VGA_BUFFER:ctrl_writedata
	wire         mm_interconnect_0_uart_avalon_jtag_slave_chipselect;               // mm_interconnect_0:UART_avalon_jtag_slave_chipselect -> UART:av_chipselect
	wire  [31:0] mm_interconnect_0_uart_avalon_jtag_slave_readdata;                 // UART:av_readdata -> mm_interconnect_0:UART_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_uart_avalon_jtag_slave_waitrequest;              // UART:av_waitrequest -> mm_interconnect_0:UART_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_uart_avalon_jtag_slave_address;                  // mm_interconnect_0:UART_avalon_jtag_slave_address -> UART:av_address
	wire         mm_interconnect_0_uart_avalon_jtag_slave_read;                     // mm_interconnect_0:UART_avalon_jtag_slave_read -> UART:av_read_n
	wire         mm_interconnect_0_uart_avalon_jtag_slave_write;                    // mm_interconnect_0:UART_avalon_jtag_slave_write -> UART:av_write_n
	wire  [31:0] mm_interconnect_0_uart_avalon_jtag_slave_writedata;                // mm_interconnect_0:UART_avalon_jtag_slave_writedata -> UART:av_writedata
	wire  [31:0] mm_interconnect_0_niosii_debug_mem_slave_readdata;                 // NIOSII:debug_mem_slave_readdata -> mm_interconnect_0:NIOSII_debug_mem_slave_readdata
	wire         mm_interconnect_0_niosii_debug_mem_slave_waitrequest;              // NIOSII:debug_mem_slave_waitrequest -> mm_interconnect_0:NIOSII_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_niosii_debug_mem_slave_debugaccess;              // mm_interconnect_0:NIOSII_debug_mem_slave_debugaccess -> NIOSII:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_niosii_debug_mem_slave_address;                  // mm_interconnect_0:NIOSII_debug_mem_slave_address -> NIOSII:debug_mem_slave_address
	wire         mm_interconnect_0_niosii_debug_mem_slave_read;                     // mm_interconnect_0:NIOSII_debug_mem_slave_read -> NIOSII:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_niosii_debug_mem_slave_byteenable;               // mm_interconnect_0:NIOSII_debug_mem_slave_byteenable -> NIOSII:debug_mem_slave_byteenable
	wire         mm_interconnect_0_niosii_debug_mem_slave_write;                    // mm_interconnect_0:NIOSII_debug_mem_slave_write -> NIOSII:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_niosii_debug_mem_slave_writedata;                // mm_interconnect_0:NIOSII_debug_mem_slave_writedata -> NIOSII:debug_mem_slave_writedata
	wire         mm_interconnect_0_timer_1s_s1_chipselect;                          // mm_interconnect_0:TIMER_1s_s1_chipselect -> TIMER_1s:chipselect
	wire  [15:0] mm_interconnect_0_timer_1s_s1_readdata;                            // TIMER_1s:readdata -> mm_interconnect_0:TIMER_1s_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_1s_s1_address;                             // mm_interconnect_0:TIMER_1s_s1_address -> TIMER_1s:address
	wire         mm_interconnect_0_timer_1s_s1_write;                               // mm_interconnect_0:TIMER_1s_s1_write -> TIMER_1s:write_n
	wire  [15:0] mm_interconnect_0_timer_1s_s1_writedata;                           // mm_interconnect_0:TIMER_1s_s1_writedata -> TIMER_1s:writedata
	wire         mm_interconnect_0_reg_7seg_s1_chipselect;                          // mm_interconnect_0:REG_7SEG_s1_chipselect -> REG_7SEG:chipselect
	wire  [31:0] mm_interconnect_0_reg_7seg_s1_readdata;                            // REG_7SEG:readdata -> mm_interconnect_0:REG_7SEG_s1_readdata
	wire   [1:0] mm_interconnect_0_reg_7seg_s1_address;                             // mm_interconnect_0:REG_7SEG_s1_address -> REG_7SEG:address
	wire         mm_interconnect_0_reg_7seg_s1_write;                               // mm_interconnect_0:REG_7SEG_s1_write -> REG_7SEG:write_n
	wire  [31:0] mm_interconnect_0_reg_7seg_s1_writedata;                           // mm_interconnect_0:REG_7SEG_s1_writedata -> REG_7SEG:writedata
	wire  [31:0] mm_interconnect_0_reg_switch_s1_readdata;                          // REG_SWITCH:readdata -> mm_interconnect_0:REG_SWITCH_s1_readdata
	wire   [1:0] mm_interconnect_0_reg_switch_s1_address;                           // mm_interconnect_0:REG_SWITCH_s1_address -> REG_SWITCH:address
	wire         mm_interconnect_0_reg_button_s1_chipselect;                        // mm_interconnect_0:REG_BUTTON_s1_chipselect -> REG_BUTTON:chipselect
	wire  [31:0] mm_interconnect_0_reg_button_s1_readdata;                          // REG_BUTTON:readdata -> mm_interconnect_0:REG_BUTTON_s1_readdata
	wire   [1:0] mm_interconnect_0_reg_button_s1_address;                           // mm_interconnect_0:REG_BUTTON_s1_address -> REG_BUTTON:address
	wire         mm_interconnect_0_reg_button_s1_write;                             // mm_interconnect_0:REG_BUTTON_s1_write -> REG_BUTTON:write_n
	wire  [31:0] mm_interconnect_0_reg_button_s1_writedata;                         // mm_interconnect_0:REG_BUTTON_s1_writedata -> REG_BUTTON:writedata
	wire         mm_interconnect_0_ram_s1_chipselect;                               // mm_interconnect_0:RAM_s1_chipselect -> RAM:chipselect
	wire  [31:0] mm_interconnect_0_ram_s1_readdata;                                 // RAM:readdata -> mm_interconnect_0:RAM_s1_readdata
	wire  [11:0] mm_interconnect_0_ram_s1_address;                                  // mm_interconnect_0:RAM_s1_address -> RAM:address
	wire   [3:0] mm_interconnect_0_ram_s1_byteenable;                               // mm_interconnect_0:RAM_s1_byteenable -> RAM:byteenable
	wire         mm_interconnect_0_ram_s1_write;                                    // mm_interconnect_0:RAM_s1_write -> RAM:write
	wire  [31:0] mm_interconnect_0_ram_s1_writedata;                                // mm_interconnect_0:RAM_s1_writedata -> RAM:writedata
	wire         mm_interconnect_0_ram_s1_clken;                                    // mm_interconnect_0:RAM_s1_clken -> RAM:clken
	wire         mm_interconnect_0_audioram_s1_chipselect;                          // mm_interconnect_0:AudioRAM_s1_chipselect -> AudioRAM:chipselect
	wire   [7:0] mm_interconnect_0_audioram_s1_readdata;                            // AudioRAM:readdata -> mm_interconnect_0:AudioRAM_s1_readdata
	wire  [14:0] mm_interconnect_0_audioram_s1_address;                             // mm_interconnect_0:AudioRAM_s1_address -> AudioRAM:address
	wire         mm_interconnect_0_audioram_s1_write;                               // mm_interconnect_0:AudioRAM_s1_write -> AudioRAM:write
	wire   [7:0] mm_interconnect_0_audioram_s1_writedata;                           // mm_interconnect_0:AudioRAM_s1_writedata -> AudioRAM:writedata
	wire         mm_interconnect_0_audioram_s1_clken;                               // mm_interconnect_0:AudioRAM_s1_clken -> AudioRAM:clken
	wire   [1:0] hps_h2f_lw_axi_master_awburst;                                     // HPS:h2f_lw_AWBURST -> mm_interconnect_1:HPS_h2f_lw_axi_master_awburst
	wire   [3:0] hps_h2f_lw_axi_master_arlen;                                       // HPS:h2f_lw_ARLEN -> mm_interconnect_1:HPS_h2f_lw_axi_master_arlen
	wire   [3:0] hps_h2f_lw_axi_master_wstrb;                                       // HPS:h2f_lw_WSTRB -> mm_interconnect_1:HPS_h2f_lw_axi_master_wstrb
	wire         hps_h2f_lw_axi_master_wready;                                      // mm_interconnect_1:HPS_h2f_lw_axi_master_wready -> HPS:h2f_lw_WREADY
	wire  [11:0] hps_h2f_lw_axi_master_rid;                                         // mm_interconnect_1:HPS_h2f_lw_axi_master_rid -> HPS:h2f_lw_RID
	wire         hps_h2f_lw_axi_master_rready;                                      // HPS:h2f_lw_RREADY -> mm_interconnect_1:HPS_h2f_lw_axi_master_rready
	wire   [3:0] hps_h2f_lw_axi_master_awlen;                                       // HPS:h2f_lw_AWLEN -> mm_interconnect_1:HPS_h2f_lw_axi_master_awlen
	wire  [11:0] hps_h2f_lw_axi_master_wid;                                         // HPS:h2f_lw_WID -> mm_interconnect_1:HPS_h2f_lw_axi_master_wid
	wire   [3:0] hps_h2f_lw_axi_master_arcache;                                     // HPS:h2f_lw_ARCACHE -> mm_interconnect_1:HPS_h2f_lw_axi_master_arcache
	wire         hps_h2f_lw_axi_master_wvalid;                                      // HPS:h2f_lw_WVALID -> mm_interconnect_1:HPS_h2f_lw_axi_master_wvalid
	wire  [20:0] hps_h2f_lw_axi_master_araddr;                                      // HPS:h2f_lw_ARADDR -> mm_interconnect_1:HPS_h2f_lw_axi_master_araddr
	wire   [2:0] hps_h2f_lw_axi_master_arprot;                                      // HPS:h2f_lw_ARPROT -> mm_interconnect_1:HPS_h2f_lw_axi_master_arprot
	wire   [2:0] hps_h2f_lw_axi_master_awprot;                                      // HPS:h2f_lw_AWPROT -> mm_interconnect_1:HPS_h2f_lw_axi_master_awprot
	wire  [31:0] hps_h2f_lw_axi_master_wdata;                                       // HPS:h2f_lw_WDATA -> mm_interconnect_1:HPS_h2f_lw_axi_master_wdata
	wire         hps_h2f_lw_axi_master_arvalid;                                     // HPS:h2f_lw_ARVALID -> mm_interconnect_1:HPS_h2f_lw_axi_master_arvalid
	wire   [3:0] hps_h2f_lw_axi_master_awcache;                                     // HPS:h2f_lw_AWCACHE -> mm_interconnect_1:HPS_h2f_lw_axi_master_awcache
	wire  [11:0] hps_h2f_lw_axi_master_arid;                                        // HPS:h2f_lw_ARID -> mm_interconnect_1:HPS_h2f_lw_axi_master_arid
	wire   [1:0] hps_h2f_lw_axi_master_arlock;                                      // HPS:h2f_lw_ARLOCK -> mm_interconnect_1:HPS_h2f_lw_axi_master_arlock
	wire   [1:0] hps_h2f_lw_axi_master_awlock;                                      // HPS:h2f_lw_AWLOCK -> mm_interconnect_1:HPS_h2f_lw_axi_master_awlock
	wire  [20:0] hps_h2f_lw_axi_master_awaddr;                                      // HPS:h2f_lw_AWADDR -> mm_interconnect_1:HPS_h2f_lw_axi_master_awaddr
	wire   [1:0] hps_h2f_lw_axi_master_bresp;                                       // mm_interconnect_1:HPS_h2f_lw_axi_master_bresp -> HPS:h2f_lw_BRESP
	wire         hps_h2f_lw_axi_master_arready;                                     // mm_interconnect_1:HPS_h2f_lw_axi_master_arready -> HPS:h2f_lw_ARREADY
	wire  [31:0] hps_h2f_lw_axi_master_rdata;                                       // mm_interconnect_1:HPS_h2f_lw_axi_master_rdata -> HPS:h2f_lw_RDATA
	wire         hps_h2f_lw_axi_master_awready;                                     // mm_interconnect_1:HPS_h2f_lw_axi_master_awready -> HPS:h2f_lw_AWREADY
	wire   [1:0] hps_h2f_lw_axi_master_arburst;                                     // HPS:h2f_lw_ARBURST -> mm_interconnect_1:HPS_h2f_lw_axi_master_arburst
	wire   [2:0] hps_h2f_lw_axi_master_arsize;                                      // HPS:h2f_lw_ARSIZE -> mm_interconnect_1:HPS_h2f_lw_axi_master_arsize
	wire         hps_h2f_lw_axi_master_bready;                                      // HPS:h2f_lw_BREADY -> mm_interconnect_1:HPS_h2f_lw_axi_master_bready
	wire         hps_h2f_lw_axi_master_rlast;                                       // mm_interconnect_1:HPS_h2f_lw_axi_master_rlast -> HPS:h2f_lw_RLAST
	wire         hps_h2f_lw_axi_master_wlast;                                       // HPS:h2f_lw_WLAST -> mm_interconnect_1:HPS_h2f_lw_axi_master_wlast
	wire   [1:0] hps_h2f_lw_axi_master_rresp;                                       // mm_interconnect_1:HPS_h2f_lw_axi_master_rresp -> HPS:h2f_lw_RRESP
	wire  [11:0] hps_h2f_lw_axi_master_awid;                                        // HPS:h2f_lw_AWID -> mm_interconnect_1:HPS_h2f_lw_axi_master_awid
	wire  [11:0] hps_h2f_lw_axi_master_bid;                                         // mm_interconnect_1:HPS_h2f_lw_axi_master_bid -> HPS:h2f_lw_BID
	wire         hps_h2f_lw_axi_master_bvalid;                                      // mm_interconnect_1:HPS_h2f_lw_axi_master_bvalid -> HPS:h2f_lw_BVALID
	wire   [2:0] hps_h2f_lw_axi_master_awsize;                                      // HPS:h2f_lw_AWSIZE -> mm_interconnect_1:HPS_h2f_lw_axi_master_awsize
	wire         hps_h2f_lw_axi_master_awvalid;                                     // HPS:h2f_lw_AWVALID -> mm_interconnect_1:HPS_h2f_lw_axi_master_awvalid
	wire         hps_h2f_lw_axi_master_rvalid;                                      // mm_interconnect_1:HPS_h2f_lw_axi_master_rvalid -> HPS:h2f_lw_RVALID
	wire         mm_interconnect_1_audioram_s2_chipselect;                          // mm_interconnect_1:AudioRAM_s2_chipselect -> AudioRAM:chipselect2
	wire   [7:0] mm_interconnect_1_audioram_s2_readdata;                            // AudioRAM:readdata2 -> mm_interconnect_1:AudioRAM_s2_readdata
	wire  [14:0] mm_interconnect_1_audioram_s2_address;                             // mm_interconnect_1:AudioRAM_s2_address -> AudioRAM:address2
	wire         mm_interconnect_1_audioram_s2_write;                               // mm_interconnect_1:AudioRAM_s2_write -> AudioRAM:write2
	wire   [7:0] mm_interconnect_1_audioram_s2_writedata;                           // mm_interconnect_1:AudioRAM_s2_writedata -> AudioRAM:writedata2
	wire         mm_interconnect_1_audioram_s2_clken;                               // mm_interconnect_1:AudioRAM_s2_clken -> AudioRAM:clken2
	wire         irq_mapper_receiver1_irq;                                          // Audio:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                          // TIMER_1s:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                          // REG_BUTTON:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                          // UART:av_irq -> irq_mapper:receiver4_irq
	wire  [31:0] niosii_irq_irq;                                                    // irq_mapper:sender_irq -> NIOSII:irq
	wire         irq_mapper_receiver0_irq;                                          // irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                                     // HPS:h2f_sdmmc_irq -> irq_synchronizer:receiver_irq
	wire         rst_controller_reset_out_reset;                                    // rst_controller:reset_out -> [Audio:reset, mm_interconnect_0:Audio_reset_reset_bridge_in_reset_reset, mm_interconnect_1:HPS_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_001_reset_out_reset;                                // rst_controller_001:reset_out -> [AudioConfig:reset, AudioRAM:reset, NIOSII:reset_n, RAM:reset, REG_7SEG:reset_n, REG_BUTTON:reset_n, REG_SWITCH:reset_n, TIMER_1s:reset_n, UART:rst_n, irq_mapper:reset, irq_synchronizer:sender_reset, mm_interconnect_0:NIOSII_reset_reset_bridge_in_reset_reset, mm_interconnect_1:AudioRAM_reset1_reset_bridge_in_reset_reset, rst_translator:in_reset]
	wire         rst_controller_001_reset_out_reset_req;                            // rst_controller_001:reset_req -> [NIOSII:reset_req, RAM:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_002_reset_out_reset;                                // rst_controller_002:reset_out -> [VGA_BUFFER:reset, VGA_CONTROLLER:reset, mm_interconnect_0:VGA_BUFFER_reset_reset_bridge_in_reset_reset]

	MP3_PC_Audio audio (
		.clk         (clk_clk),                                               //                clk.clk
		.reset       (rst_controller_reset_out_reset),                        //              reset.reset
		.address     (mm_interconnect_0_audio_avalon_audio_slave_address),    // avalon_audio_slave.address
		.chipselect  (mm_interconnect_0_audio_avalon_audio_slave_chipselect), //                   .chipselect
		.read        (mm_interconnect_0_audio_avalon_audio_slave_read),       //                   .read
		.write       (mm_interconnect_0_audio_avalon_audio_slave_write),      //                   .write
		.writedata   (mm_interconnect_0_audio_avalon_audio_slave_writedata),  //                   .writedata
		.readdata    (mm_interconnect_0_audio_avalon_audio_slave_readdata),   //                   .readdata
		.irq         (irq_mapper_receiver1_irq),                              //          interrupt.irq
		.AUD_BCLK    (audio_external_BCLK),                                   // external_interface.export
		.AUD_DACDAT  (audio_external_DACDAT),                                 //                   .export
		.AUD_DACLRCK (audio_external_DACLRCK)                                 //                   .export
	);

	MP3_PC_AudioConfig audioconfig (
		.clk         (clk_clk),                                                          //                    clk.clk
		.reset       (rst_controller_001_reset_out_reset),                               //                  reset.reset
		.address     (mm_interconnect_0_audioconfig_avalon_av_config_slave_address),     // avalon_av_config_slave.address
		.byteenable  (mm_interconnect_0_audioconfig_avalon_av_config_slave_byteenable),  //                       .byteenable
		.read        (mm_interconnect_0_audioconfig_avalon_av_config_slave_read),        //                       .read
		.write       (mm_interconnect_0_audioconfig_avalon_av_config_slave_write),       //                       .write
		.writedata   (mm_interconnect_0_audioconfig_avalon_av_config_slave_writedata),   //                       .writedata
		.readdata    (mm_interconnect_0_audioconfig_avalon_av_config_slave_readdata),    //                       .readdata
		.waitrequest (mm_interconnect_0_audioconfig_avalon_av_config_slave_waitrequest), //                       .waitrequest
		.I2C_SDAT    (audio_config_SDAT),                                                //     external_interface.export
		.I2C_SCLK    (audio_config_SCLK)                                                 //                       .export
	);

	MP3_PC_AudioPLL audiopll (
		.ref_clk_clk        (clk_clk),              //      ref_clk.clk
		.ref_reset_reset    (~hps_h2f_reset_reset), //    ref_reset.reset
		.audio_clk_clk      (audio_pll_clk_clk),    //    audio_clk.clk
		.reset_source_reset ()                      // reset_source.reset
	);

	MP3_PC_AudioRAM audioram (
		.address     (mm_interconnect_0_audioram_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_audioram_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_audioram_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_audioram_s1_write),      //       .write
		.readdata    (mm_interconnect_0_audioram_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_audioram_s1_writedata),  //       .writedata
		.address2    (mm_interconnect_1_audioram_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_1_audioram_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_1_audioram_s2_clken),      //       .clken
		.write2      (mm_interconnect_1_audioram_s2_write),      //       .write
		.readdata2   (mm_interconnect_1_audioram_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_1_audioram_s2_writedata),  //       .writedata
		.clk         (clk_clk),                                  //   clk1.clk
		.reset       (rst_controller_001_reset_out_reset),       // reset1.reset
		.freeze      (1'b0),                                     // (terminated)
		.reset_req   (1'b0)                                      // (terminated)
	);

	MP3_PC_HPS #(
		.F2S_Width (2),
		.S2F_Width (2)
	) hps (
		.h2f_mpu_eventi       (hps_h2f_mpu_events_eventi),     //      h2f_mpu_events.eventi
		.h2f_mpu_evento       (hps_h2f_mpu_events_evento),     //                    .evento
		.h2f_mpu_standbywfe   (hps_h2f_mpu_events_standbywfe), //                    .standbywfe
		.h2f_mpu_standbywfi   (hps_h2f_mpu_events_standbywfi), //                    .standbywfi
		.h2f_sdmmc_irq        (irq_synchronizer_receiver_irq), // h2f_sdmmc_interrupt.irq
		.mem_a                (memory_mem_a),                  //              memory.mem_a
		.mem_ba               (memory_mem_ba),                 //                    .mem_ba
		.mem_ck               (memory_mem_ck),                 //                    .mem_ck
		.mem_ck_n             (memory_mem_ck_n),               //                    .mem_ck_n
		.mem_cke              (memory_mem_cke),                //                    .mem_cke
		.mem_cs_n             (memory_mem_cs_n),               //                    .mem_cs_n
		.mem_ras_n            (memory_mem_ras_n),              //                    .mem_ras_n
		.mem_cas_n            (memory_mem_cas_n),              //                    .mem_cas_n
		.mem_we_n             (memory_mem_we_n),               //                    .mem_we_n
		.mem_reset_n          (memory_mem_reset_n),            //                    .mem_reset_n
		.mem_dq               (memory_mem_dq),                 //                    .mem_dq
		.mem_dqs              (memory_mem_dqs),                //                    .mem_dqs
		.mem_dqs_n            (memory_mem_dqs_n),              //                    .mem_dqs_n
		.mem_odt              (memory_mem_odt),                //                    .mem_odt
		.mem_dm               (memory_mem_dm),                 //                    .mem_dm
		.oct_rzqin            (memory_oct_rzqin),              //                    .oct_rzqin
		.hps_io_sdio_inst_CMD (hps_io_hps_io_sdio_inst_CMD),   //              hps_io.hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0  (hps_io_hps_io_sdio_inst_D0),    //                    .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1  (hps_io_hps_io_sdio_inst_D1),    //                    .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK (hps_io_hps_io_sdio_inst_CLK),   //                    .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2  (hps_io_hps_io_sdio_inst_D2),    //                    .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3  (hps_io_hps_io_sdio_inst_D3),    //                    .hps_io_sdio_inst_D3
		.h2f_rst_n            (hps_h2f_reset_reset),           //           h2f_reset.reset_n
		.f2h_sdram0_clk       (clk_clk),                       //    f2h_sdram0_clock.clk
		.f2h_sdram0_ARADDR    (),                              //     f2h_sdram0_data.araddr
		.f2h_sdram0_ARLEN     (),                              //                    .arlen
		.f2h_sdram0_ARID      (),                              //                    .arid
		.f2h_sdram0_ARSIZE    (),                              //                    .arsize
		.f2h_sdram0_ARBURST   (),                              //                    .arburst
		.f2h_sdram0_ARLOCK    (),                              //                    .arlock
		.f2h_sdram0_ARPROT    (),                              //                    .arprot
		.f2h_sdram0_ARVALID   (),                              //                    .arvalid
		.f2h_sdram0_ARCACHE   (),                              //                    .arcache
		.f2h_sdram0_AWADDR    (),                              //                    .awaddr
		.f2h_sdram0_AWLEN     (),                              //                    .awlen
		.f2h_sdram0_AWID      (),                              //                    .awid
		.f2h_sdram0_AWSIZE    (),                              //                    .awsize
		.f2h_sdram0_AWBURST   (),                              //                    .awburst
		.f2h_sdram0_AWLOCK    (),                              //                    .awlock
		.f2h_sdram0_AWPROT    (),                              //                    .awprot
		.f2h_sdram0_AWVALID   (),                              //                    .awvalid
		.f2h_sdram0_AWCACHE   (),                              //                    .awcache
		.f2h_sdram0_BRESP     (),                              //                    .bresp
		.f2h_sdram0_BID       (),                              //                    .bid
		.f2h_sdram0_BVALID    (),                              //                    .bvalid
		.f2h_sdram0_BREADY    (),                              //                    .bready
		.f2h_sdram0_ARREADY   (),                              //                    .arready
		.f2h_sdram0_AWREADY   (),                              //                    .awready
		.f2h_sdram0_RREADY    (),                              //                    .rready
		.f2h_sdram0_RDATA     (),                              //                    .rdata
		.f2h_sdram0_RRESP     (),                              //                    .rresp
		.f2h_sdram0_RLAST     (),                              //                    .rlast
		.f2h_sdram0_RID       (),                              //                    .rid
		.f2h_sdram0_RVALID    (),                              //                    .rvalid
		.f2h_sdram0_WLAST     (),                              //                    .wlast
		.f2h_sdram0_WVALID    (),                              //                    .wvalid
		.f2h_sdram0_WDATA     (),                              //                    .wdata
		.f2h_sdram0_WSTRB     (),                              //                    .wstrb
		.f2h_sdram0_WREADY    (),                              //                    .wready
		.f2h_sdram0_WID       (),                              //                    .wid
		.h2f_axi_clk          (clk_clk),                       //       h2f_axi_clock.clk
		.h2f_AWID             (),                              //      h2f_axi_master.awid
		.h2f_AWADDR           (),                              //                    .awaddr
		.h2f_AWLEN            (),                              //                    .awlen
		.h2f_AWSIZE           (),                              //                    .awsize
		.h2f_AWBURST          (),                              //                    .awburst
		.h2f_AWLOCK           (),                              //                    .awlock
		.h2f_AWCACHE          (),                              //                    .awcache
		.h2f_AWPROT           (),                              //                    .awprot
		.h2f_AWVALID          (),                              //                    .awvalid
		.h2f_AWREADY          (),                              //                    .awready
		.h2f_WID              (),                              //                    .wid
		.h2f_WDATA            (),                              //                    .wdata
		.h2f_WSTRB            (),                              //                    .wstrb
		.h2f_WLAST            (),                              //                    .wlast
		.h2f_WVALID           (),                              //                    .wvalid
		.h2f_WREADY           (),                              //                    .wready
		.h2f_BID              (),                              //                    .bid
		.h2f_BRESP            (),                              //                    .bresp
		.h2f_BVALID           (),                              //                    .bvalid
		.h2f_BREADY           (),                              //                    .bready
		.h2f_ARID             (),                              //                    .arid
		.h2f_ARADDR           (),                              //                    .araddr
		.h2f_ARLEN            (),                              //                    .arlen
		.h2f_ARSIZE           (),                              //                    .arsize
		.h2f_ARBURST          (),                              //                    .arburst
		.h2f_ARLOCK           (),                              //                    .arlock
		.h2f_ARCACHE          (),                              //                    .arcache
		.h2f_ARPROT           (),                              //                    .arprot
		.h2f_ARVALID          (),                              //                    .arvalid
		.h2f_ARREADY          (),                              //                    .arready
		.h2f_RID              (),                              //                    .rid
		.h2f_RDATA            (),                              //                    .rdata
		.h2f_RRESP            (),                              //                    .rresp
		.h2f_RLAST            (),                              //                    .rlast
		.h2f_RVALID           (),                              //                    .rvalid
		.h2f_RREADY           (),                              //                    .rready
		.f2h_axi_clk          (clk_clk),                       //       f2h_axi_clock.clk
		.f2h_AWID             (),                              //       f2h_axi_slave.awid
		.f2h_AWADDR           (),                              //                    .awaddr
		.f2h_AWLEN            (),                              //                    .awlen
		.f2h_AWSIZE           (),                              //                    .awsize
		.f2h_AWBURST          (),                              //                    .awburst
		.f2h_AWLOCK           (),                              //                    .awlock
		.f2h_AWCACHE          (),                              //                    .awcache
		.f2h_AWPROT           (),                              //                    .awprot
		.f2h_AWVALID          (),                              //                    .awvalid
		.f2h_AWREADY          (),                              //                    .awready
		.f2h_AWUSER           (),                              //                    .awuser
		.f2h_WID              (),                              //                    .wid
		.f2h_WDATA            (),                              //                    .wdata
		.f2h_WSTRB            (),                              //                    .wstrb
		.f2h_WLAST            (),                              //                    .wlast
		.f2h_WVALID           (),                              //                    .wvalid
		.f2h_WREADY           (),                              //                    .wready
		.f2h_BID              (),                              //                    .bid
		.f2h_BRESP            (),                              //                    .bresp
		.f2h_BVALID           (),                              //                    .bvalid
		.f2h_BREADY           (),                              //                    .bready
		.f2h_ARID             (),                              //                    .arid
		.f2h_ARADDR           (),                              //                    .araddr
		.f2h_ARLEN            (),                              //                    .arlen
		.f2h_ARSIZE           (),                              //                    .arsize
		.f2h_ARBURST          (),                              //                    .arburst
		.f2h_ARLOCK           (),                              //                    .arlock
		.f2h_ARCACHE          (),                              //                    .arcache
		.f2h_ARPROT           (),                              //                    .arprot
		.f2h_ARVALID          (),                              //                    .arvalid
		.f2h_ARREADY          (),                              //                    .arready
		.f2h_ARUSER           (),                              //                    .aruser
		.f2h_RID              (),                              //                    .rid
		.f2h_RDATA            (),                              //                    .rdata
		.f2h_RRESP            (),                              //                    .rresp
		.f2h_RLAST            (),                              //                    .rlast
		.f2h_RVALID           (),                              //                    .rvalid
		.f2h_RREADY           (),                              //                    .rready
		.h2f_lw_axi_clk       (clk_clk),                       //    h2f_lw_axi_clock.clk
		.h2f_lw_AWID          (hps_h2f_lw_axi_master_awid),    //   h2f_lw_axi_master.awid
		.h2f_lw_AWADDR        (hps_h2f_lw_axi_master_awaddr),  //                    .awaddr
		.h2f_lw_AWLEN         (hps_h2f_lw_axi_master_awlen),   //                    .awlen
		.h2f_lw_AWSIZE        (hps_h2f_lw_axi_master_awsize),  //                    .awsize
		.h2f_lw_AWBURST       (hps_h2f_lw_axi_master_awburst), //                    .awburst
		.h2f_lw_AWLOCK        (hps_h2f_lw_axi_master_awlock),  //                    .awlock
		.h2f_lw_AWCACHE       (hps_h2f_lw_axi_master_awcache), //                    .awcache
		.h2f_lw_AWPROT        (hps_h2f_lw_axi_master_awprot),  //                    .awprot
		.h2f_lw_AWVALID       (hps_h2f_lw_axi_master_awvalid), //                    .awvalid
		.h2f_lw_AWREADY       (hps_h2f_lw_axi_master_awready), //                    .awready
		.h2f_lw_WID           (hps_h2f_lw_axi_master_wid),     //                    .wid
		.h2f_lw_WDATA         (hps_h2f_lw_axi_master_wdata),   //                    .wdata
		.h2f_lw_WSTRB         (hps_h2f_lw_axi_master_wstrb),   //                    .wstrb
		.h2f_lw_WLAST         (hps_h2f_lw_axi_master_wlast),   //                    .wlast
		.h2f_lw_WVALID        (hps_h2f_lw_axi_master_wvalid),  //                    .wvalid
		.h2f_lw_WREADY        (hps_h2f_lw_axi_master_wready),  //                    .wready
		.h2f_lw_BID           (hps_h2f_lw_axi_master_bid),     //                    .bid
		.h2f_lw_BRESP         (hps_h2f_lw_axi_master_bresp),   //                    .bresp
		.h2f_lw_BVALID        (hps_h2f_lw_axi_master_bvalid),  //                    .bvalid
		.h2f_lw_BREADY        (hps_h2f_lw_axi_master_bready),  //                    .bready
		.h2f_lw_ARID          (hps_h2f_lw_axi_master_arid),    //                    .arid
		.h2f_lw_ARADDR        (hps_h2f_lw_axi_master_araddr),  //                    .araddr
		.h2f_lw_ARLEN         (hps_h2f_lw_axi_master_arlen),   //                    .arlen
		.h2f_lw_ARSIZE        (hps_h2f_lw_axi_master_arsize),  //                    .arsize
		.h2f_lw_ARBURST       (hps_h2f_lw_axi_master_arburst), //                    .arburst
		.h2f_lw_ARLOCK        (hps_h2f_lw_axi_master_arlock),  //                    .arlock
		.h2f_lw_ARCACHE       (hps_h2f_lw_axi_master_arcache), //                    .arcache
		.h2f_lw_ARPROT        (hps_h2f_lw_axi_master_arprot),  //                    .arprot
		.h2f_lw_ARVALID       (hps_h2f_lw_axi_master_arvalid), //                    .arvalid
		.h2f_lw_ARREADY       (hps_h2f_lw_axi_master_arready), //                    .arready
		.h2f_lw_RID           (hps_h2f_lw_axi_master_rid),     //                    .rid
		.h2f_lw_RDATA         (hps_h2f_lw_axi_master_rdata),   //                    .rdata
		.h2f_lw_RRESP         (hps_h2f_lw_axi_master_rresp),   //                    .rresp
		.h2f_lw_RLAST         (hps_h2f_lw_axi_master_rlast),   //                    .rlast
		.h2f_lw_RVALID        (hps_h2f_lw_axi_master_rvalid),  //                    .rvalid
		.h2f_lw_RREADY        (hps_h2f_lw_axi_master_rready)   //                    .rready
	);

	MP3_PC_NIOSII niosii (
		.clk                                 (clk_clk),                                              //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                  //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),               //                          .reset_req
		.d_address                           (niosii_data_master_address),                           //               data_master.address
		.d_byteenable                        (niosii_data_master_byteenable),                        //                          .byteenable
		.d_read                              (niosii_data_master_read),                              //                          .read
		.d_readdata                          (niosii_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (niosii_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (niosii_data_master_write),                             //                          .write
		.d_writedata                         (niosii_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (niosii_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (niosii_instruction_master_address),                    //        instruction_master.address
		.i_read                              (niosii_instruction_master_read),                       //                          .read
		.i_readdata                          (niosii_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (niosii_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (niosii_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (),                                                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_niosii_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_niosii_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_niosii_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_niosii_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_niosii_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_niosii_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_niosii_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_niosii_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                      // custom_instruction_master.readra
	);

	MP3_PC_PLL_VGA pll_vga (
		.refclk   (clk_clk),               //  refclk.clk
		.rst      (~hps_h2f_reset_reset),  //   reset.reset
		.outclk_0 (pll_vga_outclk0_clk),   // outclk0.clk
		.locked   (pll_vga_locked_export)  //  locked.export
	);

	MP3_PC_RAM ram (
		.clk        (clk_clk),                                //   clk1.clk
		.address    (mm_interconnect_0_ram_s1_address),       //     s1.address
		.clken      (mm_interconnect_0_ram_s1_clken),         //       .clken
		.chipselect (mm_interconnect_0_ram_s1_chipselect),    //       .chipselect
		.write      (mm_interconnect_0_ram_s1_write),         //       .write
		.readdata   (mm_interconnect_0_ram_s1_readdata),      //       .readdata
		.writedata  (mm_interconnect_0_ram_s1_writedata),     //       .writedata
		.byteenable (mm_interconnect_0_ram_s1_byteenable),    //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),     // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req), //       .reset_req
		.freeze     (1'b0)                                    // (terminated)
	);

	MP3_PC_REG_7SEG reg_7seg (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_reg_7seg_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_reg_7seg_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_reg_7seg_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_reg_7seg_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_reg_7seg_s1_readdata),   //                    .readdata
		.out_port   (seven_seg_export)                          // external_connection.export
	);

	MP3_PC_REG_BUTTON reg_button (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_reg_button_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_reg_button_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_reg_button_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_reg_button_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_reg_button_s1_readdata),   //                    .readdata
		.in_port    (buttons_export_export),                      // external_connection.export
		.irq        (irq_mapper_receiver3_irq)                    //                 irq.irq
	);

	MP3_PC_REG_SWITCH reg_switch (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_reg_switch_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_reg_switch_s1_readdata), //                    .readdata
		.in_port  (switchs_export)                            // external_connection.export
	);

	MP3_PC_TIMER_1s timer_1s (
		.clk        (clk_clk),                                  //   clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),      // reset.reset_n
		.address    (mm_interconnect_0_timer_1s_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_1s_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_1s_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_1s_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_1s_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)                  //   irq.irq
	);

	MP3_PC_UART uart (
		.clk            (clk_clk),                                              //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                  //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver4_irq)                              //               irq.irq
	);

	MP3_PC_VGA_BUFFER vga_buffer (
		.clk                  (pll_vga_outclk0_clk),                                               //                       clk.clk
		.reset                (rst_controller_002_reset_out_reset),                                //                     reset.reset
		.ctrl_address         (mm_interconnect_0_vga_buffer_avalon_char_control_slave_address),    // avalon_char_control_slave.address
		.ctrl_byteenable      (mm_interconnect_0_vga_buffer_avalon_char_control_slave_byteenable), //                          .byteenable
		.ctrl_chipselect      (mm_interconnect_0_vga_buffer_avalon_char_control_slave_chipselect), //                          .chipselect
		.ctrl_read            (mm_interconnect_0_vga_buffer_avalon_char_control_slave_read),       //                          .read
		.ctrl_write           (mm_interconnect_0_vga_buffer_avalon_char_control_slave_write),      //                          .write
		.ctrl_writedata       (mm_interconnect_0_vga_buffer_avalon_char_control_slave_writedata),  //                          .writedata
		.ctrl_readdata        (mm_interconnect_0_vga_buffer_avalon_char_control_slave_readdata),   //                          .readdata
		.buf_byteenable       (mm_interconnect_0_vga_buffer_avalon_char_buffer_slave_byteenable),  //  avalon_char_buffer_slave.byteenable
		.buf_chipselect       (mm_interconnect_0_vga_buffer_avalon_char_buffer_slave_chipselect),  //                          .chipselect
		.buf_read             (mm_interconnect_0_vga_buffer_avalon_char_buffer_slave_read),        //                          .read
		.buf_write            (mm_interconnect_0_vga_buffer_avalon_char_buffer_slave_write),       //                          .write
		.buf_writedata        (mm_interconnect_0_vga_buffer_avalon_char_buffer_slave_writedata),   //                          .writedata
		.buf_readdata         (mm_interconnect_0_vga_buffer_avalon_char_buffer_slave_readdata),    //                          .readdata
		.buf_waitrequest      (mm_interconnect_0_vga_buffer_avalon_char_buffer_slave_waitrequest), //                          .waitrequest
		.buf_address          (mm_interconnect_0_vga_buffer_avalon_char_buffer_slave_address),     //                          .address
		.stream_ready         (vga_buffer_avalon_char_source_ready),                               //        avalon_char_source.ready
		.stream_startofpacket (vga_buffer_avalon_char_source_startofpacket),                       //                          .startofpacket
		.stream_endofpacket   (vga_buffer_avalon_char_source_endofpacket),                         //                          .endofpacket
		.stream_valid         (vga_buffer_avalon_char_source_valid),                               //                          .valid
		.stream_data          (vga_buffer_avalon_char_source_data)                                 //                          .data
	);

	MP3_PC_VGA_CONTROLLER vga_controller (
		.clk           (pll_vga_outclk0_clk),                         //                clk.clk
		.reset         (rst_controller_002_reset_out_reset),          //              reset.reset
		.data          (vga_buffer_avalon_char_source_data),          //    avalon_vga_sink.data
		.startofpacket (vga_buffer_avalon_char_source_startofpacket), //                   .startofpacket
		.endofpacket   (vga_buffer_avalon_char_source_endofpacket),   //                   .endofpacket
		.valid         (vga_buffer_avalon_char_source_valid),         //                   .valid
		.ready         (vga_buffer_avalon_char_source_ready),         //                   .ready
		.VGA_CLK       (vga_controller_CLK),                          // external_interface.export
		.VGA_HS        (vga_controller_HS),                           //                   .export
		.VGA_VS        (vga_controller_VS),                           //                   .export
		.VGA_BLANK     (vga_controller_BLANK),                        //                   .export
		.VGA_SYNC      (vga_controller_SYNC),                         //                   .export
		.VGA_R         (vga_controller_R),                            //                   .export
		.VGA_G         (vga_controller_G),                            //                   .export
		.VGA_B         (vga_controller_B)                             //                   .export
	);

	MP3_PC_mm_interconnect_0 mm_interconnect_0 (
		.CLK_clk_clk                                     (clk_clk),                                                           //                                CLK_clk.clk
		.PLL_VGA_outclk0_clk                             (pll_vga_outclk0_clk),                                               //                        PLL_VGA_outclk0.clk
		.Audio_reset_reset_bridge_in_reset_reset         (rst_controller_reset_out_reset),                                    //      Audio_reset_reset_bridge_in_reset.reset
		.NIOSII_reset_reset_bridge_in_reset_reset        (rst_controller_001_reset_out_reset),                                //     NIOSII_reset_reset_bridge_in_reset.reset
		.VGA_BUFFER_reset_reset_bridge_in_reset_reset    (rst_controller_002_reset_out_reset),                                // VGA_BUFFER_reset_reset_bridge_in_reset.reset
		.NIOSII_data_master_address                      (niosii_data_master_address),                                        //                     NIOSII_data_master.address
		.NIOSII_data_master_waitrequest                  (niosii_data_master_waitrequest),                                    //                                       .waitrequest
		.NIOSII_data_master_byteenable                   (niosii_data_master_byteenable),                                     //                                       .byteenable
		.NIOSII_data_master_read                         (niosii_data_master_read),                                           //                                       .read
		.NIOSII_data_master_readdata                     (niosii_data_master_readdata),                                       //                                       .readdata
		.NIOSII_data_master_write                        (niosii_data_master_write),                                          //                                       .write
		.NIOSII_data_master_writedata                    (niosii_data_master_writedata),                                      //                                       .writedata
		.NIOSII_data_master_debugaccess                  (niosii_data_master_debugaccess),                                    //                                       .debugaccess
		.NIOSII_instruction_master_address               (niosii_instruction_master_address),                                 //              NIOSII_instruction_master.address
		.NIOSII_instruction_master_waitrequest           (niosii_instruction_master_waitrequest),                             //                                       .waitrequest
		.NIOSII_instruction_master_read                  (niosii_instruction_master_read),                                    //                                       .read
		.NIOSII_instruction_master_readdata              (niosii_instruction_master_readdata),                                //                                       .readdata
		.Audio_avalon_audio_slave_address                (mm_interconnect_0_audio_avalon_audio_slave_address),                //               Audio_avalon_audio_slave.address
		.Audio_avalon_audio_slave_write                  (mm_interconnect_0_audio_avalon_audio_slave_write),                  //                                       .write
		.Audio_avalon_audio_slave_read                   (mm_interconnect_0_audio_avalon_audio_slave_read),                   //                                       .read
		.Audio_avalon_audio_slave_readdata               (mm_interconnect_0_audio_avalon_audio_slave_readdata),               //                                       .readdata
		.Audio_avalon_audio_slave_writedata              (mm_interconnect_0_audio_avalon_audio_slave_writedata),              //                                       .writedata
		.Audio_avalon_audio_slave_chipselect             (mm_interconnect_0_audio_avalon_audio_slave_chipselect),             //                                       .chipselect
		.AudioConfig_avalon_av_config_slave_address      (mm_interconnect_0_audioconfig_avalon_av_config_slave_address),      //     AudioConfig_avalon_av_config_slave.address
		.AudioConfig_avalon_av_config_slave_write        (mm_interconnect_0_audioconfig_avalon_av_config_slave_write),        //                                       .write
		.AudioConfig_avalon_av_config_slave_read         (mm_interconnect_0_audioconfig_avalon_av_config_slave_read),         //                                       .read
		.AudioConfig_avalon_av_config_slave_readdata     (mm_interconnect_0_audioconfig_avalon_av_config_slave_readdata),     //                                       .readdata
		.AudioConfig_avalon_av_config_slave_writedata    (mm_interconnect_0_audioconfig_avalon_av_config_slave_writedata),    //                                       .writedata
		.AudioConfig_avalon_av_config_slave_byteenable   (mm_interconnect_0_audioconfig_avalon_av_config_slave_byteenable),   //                                       .byteenable
		.AudioConfig_avalon_av_config_slave_waitrequest  (mm_interconnect_0_audioconfig_avalon_av_config_slave_waitrequest),  //                                       .waitrequest
		.AudioRAM_s1_address                             (mm_interconnect_0_audioram_s1_address),                             //                            AudioRAM_s1.address
		.AudioRAM_s1_write                               (mm_interconnect_0_audioram_s1_write),                               //                                       .write
		.AudioRAM_s1_readdata                            (mm_interconnect_0_audioram_s1_readdata),                            //                                       .readdata
		.AudioRAM_s1_writedata                           (mm_interconnect_0_audioram_s1_writedata),                           //                                       .writedata
		.AudioRAM_s1_chipselect                          (mm_interconnect_0_audioram_s1_chipselect),                          //                                       .chipselect
		.AudioRAM_s1_clken                               (mm_interconnect_0_audioram_s1_clken),                               //                                       .clken
		.NIOSII_debug_mem_slave_address                  (mm_interconnect_0_niosii_debug_mem_slave_address),                  //                 NIOSII_debug_mem_slave.address
		.NIOSII_debug_mem_slave_write                    (mm_interconnect_0_niosii_debug_mem_slave_write),                    //                                       .write
		.NIOSII_debug_mem_slave_read                     (mm_interconnect_0_niosii_debug_mem_slave_read),                     //                                       .read
		.NIOSII_debug_mem_slave_readdata                 (mm_interconnect_0_niosii_debug_mem_slave_readdata),                 //                                       .readdata
		.NIOSII_debug_mem_slave_writedata                (mm_interconnect_0_niosii_debug_mem_slave_writedata),                //                                       .writedata
		.NIOSII_debug_mem_slave_byteenable               (mm_interconnect_0_niosii_debug_mem_slave_byteenable),               //                                       .byteenable
		.NIOSII_debug_mem_slave_waitrequest              (mm_interconnect_0_niosii_debug_mem_slave_waitrequest),              //                                       .waitrequest
		.NIOSII_debug_mem_slave_debugaccess              (mm_interconnect_0_niosii_debug_mem_slave_debugaccess),              //                                       .debugaccess
		.RAM_s1_address                                  (mm_interconnect_0_ram_s1_address),                                  //                                 RAM_s1.address
		.RAM_s1_write                                    (mm_interconnect_0_ram_s1_write),                                    //                                       .write
		.RAM_s1_readdata                                 (mm_interconnect_0_ram_s1_readdata),                                 //                                       .readdata
		.RAM_s1_writedata                                (mm_interconnect_0_ram_s1_writedata),                                //                                       .writedata
		.RAM_s1_byteenable                               (mm_interconnect_0_ram_s1_byteenable),                               //                                       .byteenable
		.RAM_s1_chipselect                               (mm_interconnect_0_ram_s1_chipselect),                               //                                       .chipselect
		.RAM_s1_clken                                    (mm_interconnect_0_ram_s1_clken),                                    //                                       .clken
		.REG_7SEG_s1_address                             (mm_interconnect_0_reg_7seg_s1_address),                             //                            REG_7SEG_s1.address
		.REG_7SEG_s1_write                               (mm_interconnect_0_reg_7seg_s1_write),                               //                                       .write
		.REG_7SEG_s1_readdata                            (mm_interconnect_0_reg_7seg_s1_readdata),                            //                                       .readdata
		.REG_7SEG_s1_writedata                           (mm_interconnect_0_reg_7seg_s1_writedata),                           //                                       .writedata
		.REG_7SEG_s1_chipselect                          (mm_interconnect_0_reg_7seg_s1_chipselect),                          //                                       .chipselect
		.REG_BUTTON_s1_address                           (mm_interconnect_0_reg_button_s1_address),                           //                          REG_BUTTON_s1.address
		.REG_BUTTON_s1_write                             (mm_interconnect_0_reg_button_s1_write),                             //                                       .write
		.REG_BUTTON_s1_readdata                          (mm_interconnect_0_reg_button_s1_readdata),                          //                                       .readdata
		.REG_BUTTON_s1_writedata                         (mm_interconnect_0_reg_button_s1_writedata),                         //                                       .writedata
		.REG_BUTTON_s1_chipselect                        (mm_interconnect_0_reg_button_s1_chipselect),                        //                                       .chipselect
		.REG_SWITCH_s1_address                           (mm_interconnect_0_reg_switch_s1_address),                           //                          REG_SWITCH_s1.address
		.REG_SWITCH_s1_readdata                          (mm_interconnect_0_reg_switch_s1_readdata),                          //                                       .readdata
		.TIMER_1s_s1_address                             (mm_interconnect_0_timer_1s_s1_address),                             //                            TIMER_1s_s1.address
		.TIMER_1s_s1_write                               (mm_interconnect_0_timer_1s_s1_write),                               //                                       .write
		.TIMER_1s_s1_readdata                            (mm_interconnect_0_timer_1s_s1_readdata),                            //                                       .readdata
		.TIMER_1s_s1_writedata                           (mm_interconnect_0_timer_1s_s1_writedata),                           //                                       .writedata
		.TIMER_1s_s1_chipselect                          (mm_interconnect_0_timer_1s_s1_chipselect),                          //                                       .chipselect
		.UART_avalon_jtag_slave_address                  (mm_interconnect_0_uart_avalon_jtag_slave_address),                  //                 UART_avalon_jtag_slave.address
		.UART_avalon_jtag_slave_write                    (mm_interconnect_0_uart_avalon_jtag_slave_write),                    //                                       .write
		.UART_avalon_jtag_slave_read                     (mm_interconnect_0_uart_avalon_jtag_slave_read),                     //                                       .read
		.UART_avalon_jtag_slave_readdata                 (mm_interconnect_0_uart_avalon_jtag_slave_readdata),                 //                                       .readdata
		.UART_avalon_jtag_slave_writedata                (mm_interconnect_0_uart_avalon_jtag_slave_writedata),                //                                       .writedata
		.UART_avalon_jtag_slave_waitrequest              (mm_interconnect_0_uart_avalon_jtag_slave_waitrequest),              //                                       .waitrequest
		.UART_avalon_jtag_slave_chipselect               (mm_interconnect_0_uart_avalon_jtag_slave_chipselect),               //                                       .chipselect
		.VGA_BUFFER_avalon_char_buffer_slave_address     (mm_interconnect_0_vga_buffer_avalon_char_buffer_slave_address),     //    VGA_BUFFER_avalon_char_buffer_slave.address
		.VGA_BUFFER_avalon_char_buffer_slave_write       (mm_interconnect_0_vga_buffer_avalon_char_buffer_slave_write),       //                                       .write
		.VGA_BUFFER_avalon_char_buffer_slave_read        (mm_interconnect_0_vga_buffer_avalon_char_buffer_slave_read),        //                                       .read
		.VGA_BUFFER_avalon_char_buffer_slave_readdata    (mm_interconnect_0_vga_buffer_avalon_char_buffer_slave_readdata),    //                                       .readdata
		.VGA_BUFFER_avalon_char_buffer_slave_writedata   (mm_interconnect_0_vga_buffer_avalon_char_buffer_slave_writedata),   //                                       .writedata
		.VGA_BUFFER_avalon_char_buffer_slave_byteenable  (mm_interconnect_0_vga_buffer_avalon_char_buffer_slave_byteenable),  //                                       .byteenable
		.VGA_BUFFER_avalon_char_buffer_slave_waitrequest (mm_interconnect_0_vga_buffer_avalon_char_buffer_slave_waitrequest), //                                       .waitrequest
		.VGA_BUFFER_avalon_char_buffer_slave_chipselect  (mm_interconnect_0_vga_buffer_avalon_char_buffer_slave_chipselect),  //                                       .chipselect
		.VGA_BUFFER_avalon_char_control_slave_address    (mm_interconnect_0_vga_buffer_avalon_char_control_slave_address),    //   VGA_BUFFER_avalon_char_control_slave.address
		.VGA_BUFFER_avalon_char_control_slave_write      (mm_interconnect_0_vga_buffer_avalon_char_control_slave_write),      //                                       .write
		.VGA_BUFFER_avalon_char_control_slave_read       (mm_interconnect_0_vga_buffer_avalon_char_control_slave_read),       //                                       .read
		.VGA_BUFFER_avalon_char_control_slave_readdata   (mm_interconnect_0_vga_buffer_avalon_char_control_slave_readdata),   //                                       .readdata
		.VGA_BUFFER_avalon_char_control_slave_writedata  (mm_interconnect_0_vga_buffer_avalon_char_control_slave_writedata),  //                                       .writedata
		.VGA_BUFFER_avalon_char_control_slave_byteenable (mm_interconnect_0_vga_buffer_avalon_char_control_slave_byteenable), //                                       .byteenable
		.VGA_BUFFER_avalon_char_control_slave_chipselect (mm_interconnect_0_vga_buffer_avalon_char_control_slave_chipselect)  //                                       .chipselect
	);

	MP3_PC_mm_interconnect_1 mm_interconnect_1 (
		.HPS_h2f_lw_axi_master_awid                                        (hps_h2f_lw_axi_master_awid),               //                                       HPS_h2f_lw_axi_master.awid
		.HPS_h2f_lw_axi_master_awaddr                                      (hps_h2f_lw_axi_master_awaddr),             //                                                            .awaddr
		.HPS_h2f_lw_axi_master_awlen                                       (hps_h2f_lw_axi_master_awlen),              //                                                            .awlen
		.HPS_h2f_lw_axi_master_awsize                                      (hps_h2f_lw_axi_master_awsize),             //                                                            .awsize
		.HPS_h2f_lw_axi_master_awburst                                     (hps_h2f_lw_axi_master_awburst),            //                                                            .awburst
		.HPS_h2f_lw_axi_master_awlock                                      (hps_h2f_lw_axi_master_awlock),             //                                                            .awlock
		.HPS_h2f_lw_axi_master_awcache                                     (hps_h2f_lw_axi_master_awcache),            //                                                            .awcache
		.HPS_h2f_lw_axi_master_awprot                                      (hps_h2f_lw_axi_master_awprot),             //                                                            .awprot
		.HPS_h2f_lw_axi_master_awvalid                                     (hps_h2f_lw_axi_master_awvalid),            //                                                            .awvalid
		.HPS_h2f_lw_axi_master_awready                                     (hps_h2f_lw_axi_master_awready),            //                                                            .awready
		.HPS_h2f_lw_axi_master_wid                                         (hps_h2f_lw_axi_master_wid),                //                                                            .wid
		.HPS_h2f_lw_axi_master_wdata                                       (hps_h2f_lw_axi_master_wdata),              //                                                            .wdata
		.HPS_h2f_lw_axi_master_wstrb                                       (hps_h2f_lw_axi_master_wstrb),              //                                                            .wstrb
		.HPS_h2f_lw_axi_master_wlast                                       (hps_h2f_lw_axi_master_wlast),              //                                                            .wlast
		.HPS_h2f_lw_axi_master_wvalid                                      (hps_h2f_lw_axi_master_wvalid),             //                                                            .wvalid
		.HPS_h2f_lw_axi_master_wready                                      (hps_h2f_lw_axi_master_wready),             //                                                            .wready
		.HPS_h2f_lw_axi_master_bid                                         (hps_h2f_lw_axi_master_bid),                //                                                            .bid
		.HPS_h2f_lw_axi_master_bresp                                       (hps_h2f_lw_axi_master_bresp),              //                                                            .bresp
		.HPS_h2f_lw_axi_master_bvalid                                      (hps_h2f_lw_axi_master_bvalid),             //                                                            .bvalid
		.HPS_h2f_lw_axi_master_bready                                      (hps_h2f_lw_axi_master_bready),             //                                                            .bready
		.HPS_h2f_lw_axi_master_arid                                        (hps_h2f_lw_axi_master_arid),               //                                                            .arid
		.HPS_h2f_lw_axi_master_araddr                                      (hps_h2f_lw_axi_master_araddr),             //                                                            .araddr
		.HPS_h2f_lw_axi_master_arlen                                       (hps_h2f_lw_axi_master_arlen),              //                                                            .arlen
		.HPS_h2f_lw_axi_master_arsize                                      (hps_h2f_lw_axi_master_arsize),             //                                                            .arsize
		.HPS_h2f_lw_axi_master_arburst                                     (hps_h2f_lw_axi_master_arburst),            //                                                            .arburst
		.HPS_h2f_lw_axi_master_arlock                                      (hps_h2f_lw_axi_master_arlock),             //                                                            .arlock
		.HPS_h2f_lw_axi_master_arcache                                     (hps_h2f_lw_axi_master_arcache),            //                                                            .arcache
		.HPS_h2f_lw_axi_master_arprot                                      (hps_h2f_lw_axi_master_arprot),             //                                                            .arprot
		.HPS_h2f_lw_axi_master_arvalid                                     (hps_h2f_lw_axi_master_arvalid),            //                                                            .arvalid
		.HPS_h2f_lw_axi_master_arready                                     (hps_h2f_lw_axi_master_arready),            //                                                            .arready
		.HPS_h2f_lw_axi_master_rid                                         (hps_h2f_lw_axi_master_rid),                //                                                            .rid
		.HPS_h2f_lw_axi_master_rdata                                       (hps_h2f_lw_axi_master_rdata),              //                                                            .rdata
		.HPS_h2f_lw_axi_master_rresp                                       (hps_h2f_lw_axi_master_rresp),              //                                                            .rresp
		.HPS_h2f_lw_axi_master_rlast                                       (hps_h2f_lw_axi_master_rlast),              //                                                            .rlast
		.HPS_h2f_lw_axi_master_rvalid                                      (hps_h2f_lw_axi_master_rvalid),             //                                                            .rvalid
		.HPS_h2f_lw_axi_master_rready                                      (hps_h2f_lw_axi_master_rready),             //                                                            .rready
		.CLK_clk_clk                                                       (clk_clk),                                  //                                                     CLK_clk.clk
		.AudioRAM_reset1_reset_bridge_in_reset_reset                       (rst_controller_001_reset_out_reset),       //                       AudioRAM_reset1_reset_bridge_in_reset.reset
		.HPS_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),           // HPS_h2f_lw_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.AudioRAM_s2_address                                               (mm_interconnect_1_audioram_s2_address),    //                                                 AudioRAM_s2.address
		.AudioRAM_s2_write                                                 (mm_interconnect_1_audioram_s2_write),      //                                                            .write
		.AudioRAM_s2_readdata                                              (mm_interconnect_1_audioram_s2_readdata),   //                                                            .readdata
		.AudioRAM_s2_writedata                                             (mm_interconnect_1_audioram_s2_writedata),  //                                                            .writedata
		.AudioRAM_s2_chipselect                                            (mm_interconnect_1_audioram_s2_chipselect), //                                                            .chipselect
		.AudioRAM_s2_clken                                                 (mm_interconnect_1_audioram_s2_clken)       //                                                            .clken
	);

	MP3_PC_irq_mapper irq_mapper (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),           // receiver4.irq
		.sender_irq    (niosii_irq_irq)                      //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (clk_clk),                            //       receiver_clk.clk
		.sender_clk     (clk_clk),                            //         sender_clk.clk
		.receiver_reset (),                                   // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver0_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~hps_h2f_reset_reset),           // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~hps_h2f_reset_reset),                   // reset_in0.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~hps_h2f_reset_reset),               // reset_in0.reset
		.clk            (pll_vga_outclk0_clk),                //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
